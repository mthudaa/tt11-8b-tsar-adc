magic
tech sky130A
magscale 1 2
timestamp 1746016723
<< nwell >>
rect -211 -457 211 457
<< pmos >>
rect -15 225 15 309
rect -15 47 15 131
rect -15 -131 15 -47
rect -15 -309 15 -225
<< pdiff >>
rect -73 297 -15 309
rect -73 237 -61 297
rect -27 237 -15 297
rect -73 225 -15 237
rect 15 297 73 309
rect 15 237 27 297
rect 61 237 73 297
rect 15 225 73 237
rect -73 119 -15 131
rect -73 59 -61 119
rect -27 59 -15 119
rect -73 47 -15 59
rect 15 119 73 131
rect 15 59 27 119
rect 61 59 73 119
rect 15 47 73 59
rect -73 -59 -15 -47
rect -73 -119 -61 -59
rect -27 -119 -15 -59
rect -73 -131 -15 -119
rect 15 -59 73 -47
rect 15 -119 27 -59
rect 61 -119 73 -59
rect 15 -131 73 -119
rect -73 -237 -15 -225
rect -73 -297 -61 -237
rect -27 -297 -15 -237
rect -73 -309 -15 -297
rect 15 -237 73 -225
rect 15 -297 27 -237
rect 61 -297 73 -237
rect 15 -309 73 -297
<< pdiffc >>
rect -61 237 -27 297
rect 27 237 61 297
rect -61 59 -27 119
rect 27 59 61 119
rect -61 -119 -27 -59
rect 27 -119 61 -59
rect -61 -297 -27 -237
rect 27 -297 61 -237
<< nsubdiff >>
rect -175 387 -79 421
rect 79 387 175 421
rect -175 325 -141 387
rect 141 325 175 387
rect -175 -387 -141 -325
rect 141 -387 175 -325
rect -175 -421 -79 -387
rect 79 -421 175 -387
<< nsubdiffcont >>
rect -79 387 79 421
rect -175 -325 -141 325
rect 141 -325 175 325
rect -79 -421 79 -387
<< poly >>
rect -15 309 15 335
rect -15 199 15 225
rect -15 131 15 157
rect -15 21 15 47
rect -15 -47 15 -21
rect -15 -157 15 -131
rect -15 -225 15 -199
rect -15 -335 15 -309
<< locali >>
rect -175 387 -79 421
rect 79 387 175 421
rect -175 325 -141 387
rect 141 325 175 387
rect -61 297 -27 313
rect -61 221 -27 237
rect 27 297 61 313
rect 27 221 61 237
rect -61 119 -27 135
rect -61 43 -27 59
rect 27 119 61 135
rect 27 43 61 59
rect -61 -59 -27 -43
rect -61 -135 -27 -119
rect 27 -59 61 -43
rect 27 -135 61 -119
rect -61 -237 -27 -221
rect -61 -313 -27 -297
rect 27 -237 61 -221
rect 27 -313 61 -297
rect -175 -387 -141 -325
rect 141 -387 175 -325
rect -175 -421 -79 -387
rect 79 -421 175 -387
<< viali >>
rect -61 237 -27 297
rect 27 237 61 297
rect -61 59 -27 119
rect 27 59 61 119
rect -61 -119 -27 -59
rect 27 -119 61 -59
rect -61 -297 -27 -237
rect 27 -297 61 -237
<< metal1 >>
rect -67 297 -21 309
rect -67 237 -61 297
rect -27 237 -21 297
rect -67 225 -21 237
rect 21 297 67 309
rect 21 237 27 297
rect 61 237 67 297
rect 21 225 67 237
rect -67 119 -21 131
rect -67 59 -61 119
rect -27 59 -21 119
rect -67 47 -21 59
rect 21 119 67 131
rect 21 59 27 119
rect 61 59 67 119
rect 21 47 67 59
rect -67 -59 -21 -47
rect -67 -119 -61 -59
rect -27 -119 -21 -59
rect -67 -131 -21 -119
rect 21 -59 67 -47
rect 21 -119 27 -59
rect 61 -119 67 -59
rect 21 -131 67 -119
rect -67 -237 -21 -225
rect -67 -297 -61 -237
rect -27 -297 -21 -237
rect -67 -309 -21 -297
rect 21 -237 67 -225
rect 21 -297 27 -237
rect 61 -297 67 -237
rect 21 -309 67 -297
<< properties >>
string FIXED_BBOX -158 -404 158 404
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 4 nf 1 diffcov 100 polycov 20 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
