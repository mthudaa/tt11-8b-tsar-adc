magic
tech sky130A
magscale 1 2
timestamp 1746259300
<< nwell >>
rect -246 -1439 246 1439
<< pmos >>
rect -50 920 50 1220
rect -50 492 50 792
rect -50 64 50 364
rect -50 -364 50 -64
rect -50 -792 50 -492
rect -50 -1220 50 -920
<< pdiff >>
rect -108 1208 -50 1220
rect -108 932 -96 1208
rect -62 932 -50 1208
rect -108 920 -50 932
rect 50 1208 108 1220
rect 50 932 62 1208
rect 96 932 108 1208
rect 50 920 108 932
rect -108 780 -50 792
rect -108 504 -96 780
rect -62 504 -50 780
rect -108 492 -50 504
rect 50 780 108 792
rect 50 504 62 780
rect 96 504 108 780
rect 50 492 108 504
rect -108 352 -50 364
rect -108 76 -96 352
rect -62 76 -50 352
rect -108 64 -50 76
rect 50 352 108 364
rect 50 76 62 352
rect 96 76 108 352
rect 50 64 108 76
rect -108 -76 -50 -64
rect -108 -352 -96 -76
rect -62 -352 -50 -76
rect -108 -364 -50 -352
rect 50 -76 108 -64
rect 50 -352 62 -76
rect 96 -352 108 -76
rect 50 -364 108 -352
rect -108 -504 -50 -492
rect -108 -780 -96 -504
rect -62 -780 -50 -504
rect -108 -792 -50 -780
rect 50 -504 108 -492
rect 50 -780 62 -504
rect 96 -780 108 -504
rect 50 -792 108 -780
rect -108 -932 -50 -920
rect -108 -1208 -96 -932
rect -62 -1208 -50 -932
rect -108 -1220 -50 -1208
rect 50 -932 108 -920
rect 50 -1208 62 -932
rect 96 -1208 108 -932
rect 50 -1220 108 -1208
<< pdiffc >>
rect -96 932 -62 1208
rect 62 932 96 1208
rect -96 504 -62 780
rect 62 504 96 780
rect -96 76 -62 352
rect 62 76 96 352
rect -96 -352 -62 -76
rect 62 -352 96 -76
rect -96 -780 -62 -504
rect 62 -780 96 -504
rect -96 -1208 -62 -932
rect 62 -1208 96 -932
<< nsubdiff >>
rect -210 1369 -114 1403
rect 114 1369 210 1403
rect -210 1307 -176 1369
rect 176 1307 210 1369
rect -210 -1369 -176 -1307
rect 176 -1369 210 -1307
rect -210 -1403 -114 -1369
rect 114 -1403 210 -1369
<< nsubdiffcont >>
rect -114 1369 114 1403
rect -210 -1307 -176 1307
rect 176 -1307 210 1307
rect -114 -1403 114 -1369
<< poly >>
rect -50 1301 50 1317
rect -50 1267 -34 1301
rect 34 1267 50 1301
rect -50 1220 50 1267
rect -50 873 50 920
rect -50 839 -34 873
rect 34 839 50 873
rect -50 792 50 839
rect -50 445 50 492
rect -50 411 -34 445
rect 34 411 50 445
rect -50 364 50 411
rect -50 17 50 64
rect -50 -17 -34 17
rect 34 -17 50 17
rect -50 -64 50 -17
rect -50 -411 50 -364
rect -50 -445 -34 -411
rect 34 -445 50 -411
rect -50 -492 50 -445
rect -50 -839 50 -792
rect -50 -873 -34 -839
rect 34 -873 50 -839
rect -50 -920 50 -873
rect -50 -1267 50 -1220
rect -50 -1301 -34 -1267
rect 34 -1301 50 -1267
rect -50 -1317 50 -1301
<< polycont >>
rect -34 1267 34 1301
rect -34 839 34 873
rect -34 411 34 445
rect -34 -17 34 17
rect -34 -445 34 -411
rect -34 -873 34 -839
rect -34 -1301 34 -1267
<< locali >>
rect -210 1369 -114 1403
rect 114 1369 210 1403
rect -210 1307 -176 1369
rect 176 1307 210 1369
rect -50 1267 -34 1301
rect 34 1267 50 1301
rect -96 1208 -62 1224
rect -96 916 -62 932
rect 62 1208 96 1224
rect 62 916 96 932
rect -50 839 -34 873
rect 34 839 50 873
rect -96 780 -62 796
rect -96 488 -62 504
rect 62 780 96 796
rect 62 488 96 504
rect -50 411 -34 445
rect 34 411 50 445
rect -96 352 -62 368
rect -96 60 -62 76
rect 62 352 96 368
rect 62 60 96 76
rect -50 -17 -34 17
rect 34 -17 50 17
rect -96 -76 -62 -60
rect -96 -368 -62 -352
rect 62 -76 96 -60
rect 62 -368 96 -352
rect -50 -445 -34 -411
rect 34 -445 50 -411
rect -96 -504 -62 -488
rect -96 -796 -62 -780
rect 62 -504 96 -488
rect 62 -796 96 -780
rect -50 -873 -34 -839
rect 34 -873 50 -839
rect -96 -932 -62 -916
rect -96 -1224 -62 -1208
rect 62 -932 96 -916
rect 62 -1224 96 -1208
rect -50 -1301 -34 -1267
rect 34 -1301 50 -1267
rect -210 -1369 -176 -1307
rect 176 -1369 210 -1307
rect -210 -1403 -114 -1369
rect 114 -1403 210 -1369
<< viali >>
rect -34 1267 34 1301
rect -96 932 -62 1208
rect 62 932 96 1208
rect -34 839 34 873
rect -96 504 -62 780
rect 62 504 96 780
rect -34 411 34 445
rect -96 76 -62 352
rect 62 76 96 352
rect -34 -17 34 17
rect -96 -352 -62 -76
rect 62 -352 96 -76
rect -34 -445 34 -411
rect -96 -780 -62 -504
rect 62 -780 96 -504
rect -34 -873 34 -839
rect -96 -1208 -62 -932
rect 62 -1208 96 -932
rect -34 -1301 34 -1267
<< metal1 >>
rect -46 1301 46 1307
rect -46 1267 -34 1301
rect 34 1267 46 1301
rect -46 1261 46 1267
rect -102 1208 -56 1220
rect -102 932 -96 1208
rect -62 932 -56 1208
rect -102 920 -56 932
rect 56 1208 102 1220
rect 56 932 62 1208
rect 96 932 102 1208
rect 56 920 102 932
rect -46 873 46 879
rect -46 839 -34 873
rect 34 839 46 873
rect -46 833 46 839
rect -102 780 -56 792
rect -102 504 -96 780
rect -62 504 -56 780
rect -102 492 -56 504
rect 56 780 102 792
rect 56 504 62 780
rect 96 504 102 780
rect 56 492 102 504
rect -46 445 46 451
rect -46 411 -34 445
rect 34 411 46 445
rect -46 405 46 411
rect -102 352 -56 364
rect -102 76 -96 352
rect -62 76 -56 352
rect -102 64 -56 76
rect 56 352 102 364
rect 56 76 62 352
rect 96 76 102 352
rect 56 64 102 76
rect -46 17 46 23
rect -46 -17 -34 17
rect 34 -17 46 17
rect -46 -23 46 -17
rect -102 -76 -56 -64
rect -102 -352 -96 -76
rect -62 -352 -56 -76
rect -102 -364 -56 -352
rect 56 -76 102 -64
rect 56 -352 62 -76
rect 96 -352 102 -76
rect 56 -364 102 -352
rect -46 -411 46 -405
rect -46 -445 -34 -411
rect 34 -445 46 -411
rect -46 -451 46 -445
rect -102 -504 -56 -492
rect -102 -780 -96 -504
rect -62 -780 -56 -504
rect -102 -792 -56 -780
rect 56 -504 102 -492
rect 56 -780 62 -504
rect 96 -780 102 -504
rect 56 -792 102 -780
rect -46 -839 46 -833
rect -46 -873 -34 -839
rect 34 -873 46 -839
rect -46 -879 46 -873
rect -102 -932 -56 -920
rect -102 -1208 -96 -932
rect -62 -1208 -56 -932
rect -102 -1220 -56 -1208
rect 56 -932 102 -920
rect 56 -1208 62 -932
rect 96 -1208 102 -932
rect 56 -1220 102 -1208
rect -46 -1267 46 -1261
rect -46 -1301 -34 -1267
rect 34 -1301 46 -1267
rect -46 -1307 46 -1301
<< properties >>
string FIXED_BBOX -193 -1386 193 1386
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.5 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
