magic
tech sky130A
magscale 1 2
timestamp 1746016723
<< error_p >>
rect -134 283 -76 289
rect -134 249 -122 283
rect -134 243 -76 249
rect 76 71 134 77
rect 76 37 88 71
rect 76 31 134 37
rect 76 -37 134 -31
rect 76 -71 88 -37
rect 76 -77 134 -71
rect -134 -249 -76 -243
rect -134 -283 -122 -249
rect -134 -289 -76 -283
<< nwell >>
rect -320 -421 320 421
<< pmos >>
rect -120 118 -90 202
rect 90 118 120 202
rect -120 -202 -90 -118
rect 90 -202 120 -118
<< pdiff >>
rect -182 190 -120 202
rect -182 130 -170 190
rect -136 130 -120 190
rect -182 118 -120 130
rect -90 190 -28 202
rect -90 130 -74 190
rect -40 130 -28 190
rect -90 118 -28 130
rect 28 190 90 202
rect 28 130 40 190
rect 74 130 90 190
rect 28 118 90 130
rect 120 190 182 202
rect 120 130 136 190
rect 170 130 182 190
rect 120 118 182 130
rect -182 -130 -120 -118
rect -182 -190 -170 -130
rect -136 -190 -120 -130
rect -182 -202 -120 -190
rect -90 -130 -28 -118
rect -90 -190 -74 -130
rect -40 -190 -28 -130
rect -90 -202 -28 -190
rect 28 -130 90 -118
rect 28 -190 40 -130
rect 74 -190 90 -130
rect 28 -202 90 -190
rect 120 -130 182 -118
rect 120 -190 136 -130
rect 170 -190 182 -130
rect 120 -202 182 -190
<< pdiffc >>
rect -170 130 -136 190
rect -74 130 -40 190
rect 40 130 74 190
rect 136 130 170 190
rect -170 -190 -136 -130
rect -74 -190 -40 -130
rect 40 -190 74 -130
rect 136 -190 170 -130
<< nsubdiff >>
rect -284 351 284 385
rect -284 -351 -250 351
rect 250 -351 284 351
rect -284 -385 284 -351
<< poly >>
rect -138 283 -72 299
rect -138 249 -122 283
rect -88 249 -72 283
rect -138 233 -72 249
rect -120 202 -90 233
rect 90 202 120 228
rect -120 92 -90 118
rect 90 87 120 118
rect 72 71 138 87
rect 72 37 88 71
rect 122 37 138 71
rect 72 21 138 37
rect 72 -37 138 -21
rect 72 -71 88 -37
rect 122 -71 138 -37
rect 72 -87 138 -71
rect -120 -118 -90 -92
rect 90 -118 120 -87
rect -120 -233 -90 -202
rect 90 -228 120 -202
rect -138 -249 -72 -233
rect -138 -283 -122 -249
rect -88 -283 -72 -249
rect -138 -299 -72 -283
<< polycont >>
rect -122 249 -88 283
rect 88 37 122 71
rect 88 -71 122 -37
rect -122 -283 -88 -249
<< locali >>
rect -138 249 -122 283
rect -88 249 -72 283
rect -170 190 -136 206
rect -170 114 -136 130
rect -74 190 -40 206
rect -74 114 -40 130
rect 40 190 74 206
rect 40 114 74 130
rect 136 190 170 206
rect 136 114 170 130
rect 72 37 88 71
rect 122 37 138 71
rect 72 -71 88 -37
rect 122 -71 138 -37
rect -170 -130 -136 -114
rect -170 -206 -136 -190
rect -74 -130 -40 -114
rect -74 -206 -40 -190
rect 40 -130 74 -114
rect 40 -206 74 -190
rect 136 -130 170 -114
rect 136 -206 170 -190
rect -138 -283 -122 -249
rect -88 -283 -72 -249
<< viali >>
rect -122 249 -88 283
rect -170 130 -136 190
rect -74 130 -40 190
rect 40 130 74 190
rect 136 130 170 190
rect 88 37 122 71
rect 88 -71 122 -37
rect -170 -190 -136 -130
rect -74 -190 -40 -130
rect 40 -190 74 -130
rect 136 -190 170 -130
rect -122 -283 -88 -249
<< metal1 >>
rect -134 283 -76 289
rect -134 249 -122 283
rect -88 249 -76 283
rect -134 243 -76 249
rect -176 190 -130 202
rect -176 130 -170 190
rect -136 130 -130 190
rect -176 118 -130 130
rect -80 190 -34 202
rect -80 130 -74 190
rect -40 130 -34 190
rect -80 118 -34 130
rect 34 190 80 202
rect 34 130 40 190
rect 74 130 80 190
rect 34 118 80 130
rect 130 190 176 202
rect 130 130 136 190
rect 170 130 176 190
rect 130 118 176 130
rect 76 71 134 77
rect 76 37 88 71
rect 122 37 134 71
rect 76 31 134 37
rect 76 -37 134 -31
rect 76 -71 88 -37
rect 122 -71 134 -37
rect 76 -77 134 -71
rect -176 -130 -130 -118
rect -176 -190 -170 -130
rect -136 -190 -130 -130
rect -176 -202 -130 -190
rect -80 -130 -34 -118
rect -80 -190 -74 -130
rect -40 -190 -34 -130
rect -80 -202 -34 -190
rect 34 -130 80 -118
rect 34 -190 40 -130
rect 74 -190 80 -130
rect 34 -202 80 -190
rect 130 -130 176 -118
rect 130 -190 136 -130
rect 170 -190 176 -130
rect 130 -202 176 -190
rect -134 -249 -76 -243
rect -134 -283 -122 -249
rect -88 -283 -76 -249
rect -134 -289 -76 -283
<< properties >>
string FIXED_BBOX -267 -368 267 368
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 2 nf 2 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
