magic
tech sky130A
magscale 1 2
timestamp 1746259300
<< pwell >>
rect -246 -785 246 785
<< nmos >>
rect -50 475 50 575
rect -50 265 50 365
rect -50 55 50 155
rect -50 -155 50 -55
rect -50 -365 50 -265
rect -50 -575 50 -475
<< ndiff >>
rect -108 563 -50 575
rect -108 487 -96 563
rect -62 487 -50 563
rect -108 475 -50 487
rect 50 563 108 575
rect 50 487 62 563
rect 96 487 108 563
rect 50 475 108 487
rect -108 353 -50 365
rect -108 277 -96 353
rect -62 277 -50 353
rect -108 265 -50 277
rect 50 353 108 365
rect 50 277 62 353
rect 96 277 108 353
rect 50 265 108 277
rect -108 143 -50 155
rect -108 67 -96 143
rect -62 67 -50 143
rect -108 55 -50 67
rect 50 143 108 155
rect 50 67 62 143
rect 96 67 108 143
rect 50 55 108 67
rect -108 -67 -50 -55
rect -108 -143 -96 -67
rect -62 -143 -50 -67
rect -108 -155 -50 -143
rect 50 -67 108 -55
rect 50 -143 62 -67
rect 96 -143 108 -67
rect 50 -155 108 -143
rect -108 -277 -50 -265
rect -108 -353 -96 -277
rect -62 -353 -50 -277
rect -108 -365 -50 -353
rect 50 -277 108 -265
rect 50 -353 62 -277
rect 96 -353 108 -277
rect 50 -365 108 -353
rect -108 -487 -50 -475
rect -108 -563 -96 -487
rect -62 -563 -50 -487
rect -108 -575 -50 -563
rect 50 -487 108 -475
rect 50 -563 62 -487
rect 96 -563 108 -487
rect 50 -575 108 -563
<< ndiffc >>
rect -96 487 -62 563
rect 62 487 96 563
rect -96 277 -62 353
rect 62 277 96 353
rect -96 67 -62 143
rect 62 67 96 143
rect -96 -143 -62 -67
rect 62 -143 96 -67
rect -96 -353 -62 -277
rect 62 -353 96 -277
rect -96 -563 -62 -487
rect 62 -563 96 -487
<< psubdiff >>
rect -210 715 -114 749
rect 114 715 210 749
rect -210 653 -176 715
rect 176 653 210 715
rect -210 -715 -176 -653
rect 176 -715 210 -653
rect -210 -749 -114 -715
rect 114 -749 210 -715
<< psubdiffcont >>
rect -114 715 114 749
rect -210 -653 -176 653
rect 176 -653 210 653
rect -114 -749 114 -715
<< poly >>
rect -50 647 50 663
rect -50 613 -34 647
rect 34 613 50 647
rect -50 575 50 613
rect -50 437 50 475
rect -50 403 -34 437
rect 34 403 50 437
rect -50 365 50 403
rect -50 227 50 265
rect -50 193 -34 227
rect 34 193 50 227
rect -50 155 50 193
rect -50 17 50 55
rect -50 -17 -34 17
rect 34 -17 50 17
rect -50 -55 50 -17
rect -50 -193 50 -155
rect -50 -227 -34 -193
rect 34 -227 50 -193
rect -50 -265 50 -227
rect -50 -403 50 -365
rect -50 -437 -34 -403
rect 34 -437 50 -403
rect -50 -475 50 -437
rect -50 -613 50 -575
rect -50 -647 -34 -613
rect 34 -647 50 -613
rect -50 -663 50 -647
<< polycont >>
rect -34 613 34 647
rect -34 403 34 437
rect -34 193 34 227
rect -34 -17 34 17
rect -34 -227 34 -193
rect -34 -437 34 -403
rect -34 -647 34 -613
<< locali >>
rect -210 715 -114 749
rect 114 715 210 749
rect -210 653 -176 715
rect 176 653 210 715
rect -50 613 -34 647
rect 34 613 50 647
rect -96 563 -62 579
rect -96 471 -62 487
rect 62 563 96 579
rect 62 471 96 487
rect -50 403 -34 437
rect 34 403 50 437
rect -96 353 -62 369
rect -96 261 -62 277
rect 62 353 96 369
rect 62 261 96 277
rect -50 193 -34 227
rect 34 193 50 227
rect -96 143 -62 159
rect -96 51 -62 67
rect 62 143 96 159
rect 62 51 96 67
rect -50 -17 -34 17
rect 34 -17 50 17
rect -96 -67 -62 -51
rect -96 -159 -62 -143
rect 62 -67 96 -51
rect 62 -159 96 -143
rect -50 -227 -34 -193
rect 34 -227 50 -193
rect -96 -277 -62 -261
rect -96 -369 -62 -353
rect 62 -277 96 -261
rect 62 -369 96 -353
rect -50 -437 -34 -403
rect 34 -437 50 -403
rect -96 -487 -62 -471
rect -96 -579 -62 -563
rect 62 -487 96 -471
rect 62 -579 96 -563
rect -50 -647 -34 -613
rect 34 -647 50 -613
rect -210 -715 -176 -653
rect 176 -715 210 -653
rect -210 -749 -114 -715
rect 114 -749 210 -715
<< viali >>
rect -34 613 34 647
rect -96 487 -62 563
rect 62 487 96 563
rect -34 403 34 437
rect -96 277 -62 353
rect 62 277 96 353
rect -34 193 34 227
rect -96 67 -62 143
rect 62 67 96 143
rect -34 -17 34 17
rect -96 -143 -62 -67
rect 62 -143 96 -67
rect -34 -227 34 -193
rect -96 -353 -62 -277
rect 62 -353 96 -277
rect -34 -437 34 -403
rect -96 -563 -62 -487
rect 62 -563 96 -487
rect -34 -647 34 -613
<< metal1 >>
rect -46 647 46 653
rect -46 613 -34 647
rect 34 613 46 647
rect -46 607 46 613
rect -102 563 -56 575
rect -102 487 -96 563
rect -62 487 -56 563
rect -102 475 -56 487
rect 56 563 102 575
rect 56 487 62 563
rect 96 487 102 563
rect 56 475 102 487
rect -46 437 46 443
rect -46 403 -34 437
rect 34 403 46 437
rect -46 397 46 403
rect -102 353 -56 365
rect -102 277 -96 353
rect -62 277 -56 353
rect -102 265 -56 277
rect 56 353 102 365
rect 56 277 62 353
rect 96 277 102 353
rect 56 265 102 277
rect -46 227 46 233
rect -46 193 -34 227
rect 34 193 46 227
rect -46 187 46 193
rect -102 143 -56 155
rect -102 67 -96 143
rect -62 67 -56 143
rect -102 55 -56 67
rect 56 143 102 155
rect 56 67 62 143
rect 96 67 102 143
rect 56 55 102 67
rect -46 17 46 23
rect -46 -17 -34 17
rect 34 -17 46 17
rect -46 -23 46 -17
rect -102 -67 -56 -55
rect -102 -143 -96 -67
rect -62 -143 -56 -67
rect -102 -155 -56 -143
rect 56 -67 102 -55
rect 56 -143 62 -67
rect 96 -143 102 -67
rect 56 -155 102 -143
rect -46 -193 46 -187
rect -46 -227 -34 -193
rect 34 -227 46 -193
rect -46 -233 46 -227
rect -102 -277 -56 -265
rect -102 -353 -96 -277
rect -62 -353 -56 -277
rect -102 -365 -56 -353
rect 56 -277 102 -265
rect 56 -353 62 -277
rect 96 -353 102 -277
rect 56 -365 102 -353
rect -46 -403 46 -397
rect -46 -437 -34 -403
rect 34 -437 46 -403
rect -46 -443 46 -437
rect -102 -487 -56 -475
rect -102 -563 -96 -487
rect -62 -563 -56 -487
rect -102 -575 -56 -563
rect 56 -487 102 -475
rect 56 -563 62 -487
rect 96 -563 102 -487
rect 56 -575 102 -563
rect -46 -613 46 -607
rect -46 -647 -34 -613
rect 34 -647 46 -613
rect -46 -653 46 -647
<< properties >>
string FIXED_BBOX -193 -732 193 732
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.5 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
