magic
tech sky130A
magscale 1 2
timestamp 1747688232
<< metal3 >>
rect -23884 18892 -22712 18920
rect -23884 18068 -22796 18892
rect -22732 18068 -22712 18892
rect -23884 18040 -22712 18068
rect -22472 18892 -21300 18920
rect -22472 18068 -21384 18892
rect -21320 18068 -21300 18892
rect -22472 18040 -21300 18068
rect -21060 18892 -19888 18920
rect -21060 18068 -19972 18892
rect -19908 18068 -19888 18892
rect -21060 18040 -19888 18068
rect -19648 18892 -18476 18920
rect -19648 18068 -18560 18892
rect -18496 18068 -18476 18892
rect -19648 18040 -18476 18068
rect -18236 18892 -17064 18920
rect -18236 18068 -17148 18892
rect -17084 18068 -17064 18892
rect -18236 18040 -17064 18068
rect -16824 18892 -15652 18920
rect -16824 18068 -15736 18892
rect -15672 18068 -15652 18892
rect -16824 18040 -15652 18068
rect -15412 18892 -14240 18920
rect -15412 18068 -14324 18892
rect -14260 18068 -14240 18892
rect -15412 18040 -14240 18068
rect -14000 18892 -12828 18920
rect -14000 18068 -12912 18892
rect -12848 18068 -12828 18892
rect -14000 18040 -12828 18068
rect -12588 18892 -11416 18920
rect -12588 18068 -11500 18892
rect -11436 18068 -11416 18892
rect -12588 18040 -11416 18068
rect -11176 18892 -10004 18920
rect -11176 18068 -10088 18892
rect -10024 18068 -10004 18892
rect -11176 18040 -10004 18068
rect -9764 18892 -8592 18920
rect -9764 18068 -8676 18892
rect -8612 18068 -8592 18892
rect -9764 18040 -8592 18068
rect -8352 18892 -7180 18920
rect -8352 18068 -7264 18892
rect -7200 18068 -7180 18892
rect -8352 18040 -7180 18068
rect -6940 18892 -5768 18920
rect -6940 18068 -5852 18892
rect -5788 18068 -5768 18892
rect -6940 18040 -5768 18068
rect -5528 18892 -4356 18920
rect -5528 18068 -4440 18892
rect -4376 18068 -4356 18892
rect -5528 18040 -4356 18068
rect -4116 18892 -2944 18920
rect -4116 18068 -3028 18892
rect -2964 18068 -2944 18892
rect -4116 18040 -2944 18068
rect -2704 18892 -1532 18920
rect -2704 18068 -1616 18892
rect -1552 18068 -1532 18892
rect -2704 18040 -1532 18068
rect -1292 18892 -120 18920
rect -1292 18068 -204 18892
rect -140 18068 -120 18892
rect -1292 18040 -120 18068
rect 120 18892 1292 18920
rect 120 18068 1208 18892
rect 1272 18068 1292 18892
rect 120 18040 1292 18068
rect 1532 18892 2704 18920
rect 1532 18068 2620 18892
rect 2684 18068 2704 18892
rect 1532 18040 2704 18068
rect 2944 18892 4116 18920
rect 2944 18068 4032 18892
rect 4096 18068 4116 18892
rect 2944 18040 4116 18068
rect 4356 18892 5528 18920
rect 4356 18068 5444 18892
rect 5508 18068 5528 18892
rect 4356 18040 5528 18068
rect 5768 18892 6940 18920
rect 5768 18068 6856 18892
rect 6920 18068 6940 18892
rect 5768 18040 6940 18068
rect 7180 18892 8352 18920
rect 7180 18068 8268 18892
rect 8332 18068 8352 18892
rect 7180 18040 8352 18068
rect 8592 18892 9764 18920
rect 8592 18068 9680 18892
rect 9744 18068 9764 18892
rect 8592 18040 9764 18068
rect 10004 18892 11176 18920
rect 10004 18068 11092 18892
rect 11156 18068 11176 18892
rect 10004 18040 11176 18068
rect 11416 18892 12588 18920
rect 11416 18068 12504 18892
rect 12568 18068 12588 18892
rect 11416 18040 12588 18068
rect 12828 18892 14000 18920
rect 12828 18068 13916 18892
rect 13980 18068 14000 18892
rect 12828 18040 14000 18068
rect 14240 18892 15412 18920
rect 14240 18068 15328 18892
rect 15392 18068 15412 18892
rect 14240 18040 15412 18068
rect 15652 18892 16824 18920
rect 15652 18068 16740 18892
rect 16804 18068 16824 18892
rect 15652 18040 16824 18068
rect 17064 18892 18236 18920
rect 17064 18068 18152 18892
rect 18216 18068 18236 18892
rect 17064 18040 18236 18068
rect 18476 18892 19648 18920
rect 18476 18068 19564 18892
rect 19628 18068 19648 18892
rect 18476 18040 19648 18068
rect 19888 18892 21060 18920
rect 19888 18068 20976 18892
rect 21040 18068 21060 18892
rect 19888 18040 21060 18068
rect 21300 18892 22472 18920
rect 21300 18068 22388 18892
rect 22452 18068 22472 18892
rect 21300 18040 22472 18068
rect 22712 18892 23884 18920
rect 22712 18068 23800 18892
rect 23864 18068 23884 18892
rect 22712 18040 23884 18068
rect -23884 17772 -22712 17800
rect -23884 16948 -22796 17772
rect -22732 16948 -22712 17772
rect -23884 16920 -22712 16948
rect -22472 17772 -21300 17800
rect -22472 16948 -21384 17772
rect -21320 16948 -21300 17772
rect -22472 16920 -21300 16948
rect -21060 17772 -19888 17800
rect -21060 16948 -19972 17772
rect -19908 16948 -19888 17772
rect -21060 16920 -19888 16948
rect -19648 17772 -18476 17800
rect -19648 16948 -18560 17772
rect -18496 16948 -18476 17772
rect -19648 16920 -18476 16948
rect -18236 17772 -17064 17800
rect -18236 16948 -17148 17772
rect -17084 16948 -17064 17772
rect -18236 16920 -17064 16948
rect -16824 17772 -15652 17800
rect -16824 16948 -15736 17772
rect -15672 16948 -15652 17772
rect -16824 16920 -15652 16948
rect -15412 17772 -14240 17800
rect -15412 16948 -14324 17772
rect -14260 16948 -14240 17772
rect -15412 16920 -14240 16948
rect -14000 17772 -12828 17800
rect -14000 16948 -12912 17772
rect -12848 16948 -12828 17772
rect -14000 16920 -12828 16948
rect -12588 17772 -11416 17800
rect -12588 16948 -11500 17772
rect -11436 16948 -11416 17772
rect -12588 16920 -11416 16948
rect -11176 17772 -10004 17800
rect -11176 16948 -10088 17772
rect -10024 16948 -10004 17772
rect -11176 16920 -10004 16948
rect -9764 17772 -8592 17800
rect -9764 16948 -8676 17772
rect -8612 16948 -8592 17772
rect -9764 16920 -8592 16948
rect -8352 17772 -7180 17800
rect -8352 16948 -7264 17772
rect -7200 16948 -7180 17772
rect -8352 16920 -7180 16948
rect -6940 17772 -5768 17800
rect -6940 16948 -5852 17772
rect -5788 16948 -5768 17772
rect -6940 16920 -5768 16948
rect -5528 17772 -4356 17800
rect -5528 16948 -4440 17772
rect -4376 16948 -4356 17772
rect -5528 16920 -4356 16948
rect -4116 17772 -2944 17800
rect -4116 16948 -3028 17772
rect -2964 16948 -2944 17772
rect -4116 16920 -2944 16948
rect -2704 17772 -1532 17800
rect -2704 16948 -1616 17772
rect -1552 16948 -1532 17772
rect -2704 16920 -1532 16948
rect -1292 17772 -120 17800
rect -1292 16948 -204 17772
rect -140 16948 -120 17772
rect -1292 16920 -120 16948
rect 120 17772 1292 17800
rect 120 16948 1208 17772
rect 1272 16948 1292 17772
rect 120 16920 1292 16948
rect 1532 17772 2704 17800
rect 1532 16948 2620 17772
rect 2684 16948 2704 17772
rect 1532 16920 2704 16948
rect 2944 17772 4116 17800
rect 2944 16948 4032 17772
rect 4096 16948 4116 17772
rect 2944 16920 4116 16948
rect 4356 17772 5528 17800
rect 4356 16948 5444 17772
rect 5508 16948 5528 17772
rect 4356 16920 5528 16948
rect 5768 17772 6940 17800
rect 5768 16948 6856 17772
rect 6920 16948 6940 17772
rect 5768 16920 6940 16948
rect 7180 17772 8352 17800
rect 7180 16948 8268 17772
rect 8332 16948 8352 17772
rect 7180 16920 8352 16948
rect 8592 17772 9764 17800
rect 8592 16948 9680 17772
rect 9744 16948 9764 17772
rect 8592 16920 9764 16948
rect 10004 17772 11176 17800
rect 10004 16948 11092 17772
rect 11156 16948 11176 17772
rect 10004 16920 11176 16948
rect 11416 17772 12588 17800
rect 11416 16948 12504 17772
rect 12568 16948 12588 17772
rect 11416 16920 12588 16948
rect 12828 17772 14000 17800
rect 12828 16948 13916 17772
rect 13980 16948 14000 17772
rect 12828 16920 14000 16948
rect 14240 17772 15412 17800
rect 14240 16948 15328 17772
rect 15392 16948 15412 17772
rect 14240 16920 15412 16948
rect 15652 17772 16824 17800
rect 15652 16948 16740 17772
rect 16804 16948 16824 17772
rect 15652 16920 16824 16948
rect 17064 17772 18236 17800
rect 17064 16948 18152 17772
rect 18216 16948 18236 17772
rect 17064 16920 18236 16948
rect 18476 17772 19648 17800
rect 18476 16948 19564 17772
rect 19628 16948 19648 17772
rect 18476 16920 19648 16948
rect 19888 17772 21060 17800
rect 19888 16948 20976 17772
rect 21040 16948 21060 17772
rect 19888 16920 21060 16948
rect 21300 17772 22472 17800
rect 21300 16948 22388 17772
rect 22452 16948 22472 17772
rect 21300 16920 22472 16948
rect 22712 17772 23884 17800
rect 22712 16948 23800 17772
rect 23864 16948 23884 17772
rect 22712 16920 23884 16948
rect -23884 16652 -22712 16680
rect -23884 15828 -22796 16652
rect -22732 15828 -22712 16652
rect -23884 15800 -22712 15828
rect -22472 16652 -21300 16680
rect -22472 15828 -21384 16652
rect -21320 15828 -21300 16652
rect -22472 15800 -21300 15828
rect -21060 16652 -19888 16680
rect -21060 15828 -19972 16652
rect -19908 15828 -19888 16652
rect -21060 15800 -19888 15828
rect -19648 16652 -18476 16680
rect -19648 15828 -18560 16652
rect -18496 15828 -18476 16652
rect -19648 15800 -18476 15828
rect -18236 16652 -17064 16680
rect -18236 15828 -17148 16652
rect -17084 15828 -17064 16652
rect -18236 15800 -17064 15828
rect -16824 16652 -15652 16680
rect -16824 15828 -15736 16652
rect -15672 15828 -15652 16652
rect -16824 15800 -15652 15828
rect -15412 16652 -14240 16680
rect -15412 15828 -14324 16652
rect -14260 15828 -14240 16652
rect -15412 15800 -14240 15828
rect -14000 16652 -12828 16680
rect -14000 15828 -12912 16652
rect -12848 15828 -12828 16652
rect -14000 15800 -12828 15828
rect -12588 16652 -11416 16680
rect -12588 15828 -11500 16652
rect -11436 15828 -11416 16652
rect -12588 15800 -11416 15828
rect -11176 16652 -10004 16680
rect -11176 15828 -10088 16652
rect -10024 15828 -10004 16652
rect -11176 15800 -10004 15828
rect -9764 16652 -8592 16680
rect -9764 15828 -8676 16652
rect -8612 15828 -8592 16652
rect -9764 15800 -8592 15828
rect -8352 16652 -7180 16680
rect -8352 15828 -7264 16652
rect -7200 15828 -7180 16652
rect -8352 15800 -7180 15828
rect -6940 16652 -5768 16680
rect -6940 15828 -5852 16652
rect -5788 15828 -5768 16652
rect -6940 15800 -5768 15828
rect -5528 16652 -4356 16680
rect -5528 15828 -4440 16652
rect -4376 15828 -4356 16652
rect -5528 15800 -4356 15828
rect -4116 16652 -2944 16680
rect -4116 15828 -3028 16652
rect -2964 15828 -2944 16652
rect -4116 15800 -2944 15828
rect -2704 16652 -1532 16680
rect -2704 15828 -1616 16652
rect -1552 15828 -1532 16652
rect -2704 15800 -1532 15828
rect -1292 16652 -120 16680
rect -1292 15828 -204 16652
rect -140 15828 -120 16652
rect -1292 15800 -120 15828
rect 120 16652 1292 16680
rect 120 15828 1208 16652
rect 1272 15828 1292 16652
rect 120 15800 1292 15828
rect 1532 16652 2704 16680
rect 1532 15828 2620 16652
rect 2684 15828 2704 16652
rect 1532 15800 2704 15828
rect 2944 16652 4116 16680
rect 2944 15828 4032 16652
rect 4096 15828 4116 16652
rect 2944 15800 4116 15828
rect 4356 16652 5528 16680
rect 4356 15828 5444 16652
rect 5508 15828 5528 16652
rect 4356 15800 5528 15828
rect 5768 16652 6940 16680
rect 5768 15828 6856 16652
rect 6920 15828 6940 16652
rect 5768 15800 6940 15828
rect 7180 16652 8352 16680
rect 7180 15828 8268 16652
rect 8332 15828 8352 16652
rect 7180 15800 8352 15828
rect 8592 16652 9764 16680
rect 8592 15828 9680 16652
rect 9744 15828 9764 16652
rect 8592 15800 9764 15828
rect 10004 16652 11176 16680
rect 10004 15828 11092 16652
rect 11156 15828 11176 16652
rect 10004 15800 11176 15828
rect 11416 16652 12588 16680
rect 11416 15828 12504 16652
rect 12568 15828 12588 16652
rect 11416 15800 12588 15828
rect 12828 16652 14000 16680
rect 12828 15828 13916 16652
rect 13980 15828 14000 16652
rect 12828 15800 14000 15828
rect 14240 16652 15412 16680
rect 14240 15828 15328 16652
rect 15392 15828 15412 16652
rect 14240 15800 15412 15828
rect 15652 16652 16824 16680
rect 15652 15828 16740 16652
rect 16804 15828 16824 16652
rect 15652 15800 16824 15828
rect 17064 16652 18236 16680
rect 17064 15828 18152 16652
rect 18216 15828 18236 16652
rect 17064 15800 18236 15828
rect 18476 16652 19648 16680
rect 18476 15828 19564 16652
rect 19628 15828 19648 16652
rect 18476 15800 19648 15828
rect 19888 16652 21060 16680
rect 19888 15828 20976 16652
rect 21040 15828 21060 16652
rect 19888 15800 21060 15828
rect 21300 16652 22472 16680
rect 21300 15828 22388 16652
rect 22452 15828 22472 16652
rect 21300 15800 22472 15828
rect 22712 16652 23884 16680
rect 22712 15828 23800 16652
rect 23864 15828 23884 16652
rect 22712 15800 23884 15828
rect -23884 15532 -22712 15560
rect -23884 14708 -22796 15532
rect -22732 14708 -22712 15532
rect -23884 14680 -22712 14708
rect -22472 15532 -21300 15560
rect -22472 14708 -21384 15532
rect -21320 14708 -21300 15532
rect -22472 14680 -21300 14708
rect -21060 15532 -19888 15560
rect -21060 14708 -19972 15532
rect -19908 14708 -19888 15532
rect -21060 14680 -19888 14708
rect -19648 15532 -18476 15560
rect -19648 14708 -18560 15532
rect -18496 14708 -18476 15532
rect -19648 14680 -18476 14708
rect -18236 15532 -17064 15560
rect -18236 14708 -17148 15532
rect -17084 14708 -17064 15532
rect -18236 14680 -17064 14708
rect -16824 15532 -15652 15560
rect -16824 14708 -15736 15532
rect -15672 14708 -15652 15532
rect -16824 14680 -15652 14708
rect -15412 15532 -14240 15560
rect -15412 14708 -14324 15532
rect -14260 14708 -14240 15532
rect -15412 14680 -14240 14708
rect -14000 15532 -12828 15560
rect -14000 14708 -12912 15532
rect -12848 14708 -12828 15532
rect -14000 14680 -12828 14708
rect -12588 15532 -11416 15560
rect -12588 14708 -11500 15532
rect -11436 14708 -11416 15532
rect -12588 14680 -11416 14708
rect -11176 15532 -10004 15560
rect -11176 14708 -10088 15532
rect -10024 14708 -10004 15532
rect -11176 14680 -10004 14708
rect -9764 15532 -8592 15560
rect -9764 14708 -8676 15532
rect -8612 14708 -8592 15532
rect -9764 14680 -8592 14708
rect -8352 15532 -7180 15560
rect -8352 14708 -7264 15532
rect -7200 14708 -7180 15532
rect -8352 14680 -7180 14708
rect -6940 15532 -5768 15560
rect -6940 14708 -5852 15532
rect -5788 14708 -5768 15532
rect -6940 14680 -5768 14708
rect -5528 15532 -4356 15560
rect -5528 14708 -4440 15532
rect -4376 14708 -4356 15532
rect -5528 14680 -4356 14708
rect -4116 15532 -2944 15560
rect -4116 14708 -3028 15532
rect -2964 14708 -2944 15532
rect -4116 14680 -2944 14708
rect -2704 15532 -1532 15560
rect -2704 14708 -1616 15532
rect -1552 14708 -1532 15532
rect -2704 14680 -1532 14708
rect -1292 15532 -120 15560
rect -1292 14708 -204 15532
rect -140 14708 -120 15532
rect -1292 14680 -120 14708
rect 120 15532 1292 15560
rect 120 14708 1208 15532
rect 1272 14708 1292 15532
rect 120 14680 1292 14708
rect 1532 15532 2704 15560
rect 1532 14708 2620 15532
rect 2684 14708 2704 15532
rect 1532 14680 2704 14708
rect 2944 15532 4116 15560
rect 2944 14708 4032 15532
rect 4096 14708 4116 15532
rect 2944 14680 4116 14708
rect 4356 15532 5528 15560
rect 4356 14708 5444 15532
rect 5508 14708 5528 15532
rect 4356 14680 5528 14708
rect 5768 15532 6940 15560
rect 5768 14708 6856 15532
rect 6920 14708 6940 15532
rect 5768 14680 6940 14708
rect 7180 15532 8352 15560
rect 7180 14708 8268 15532
rect 8332 14708 8352 15532
rect 7180 14680 8352 14708
rect 8592 15532 9764 15560
rect 8592 14708 9680 15532
rect 9744 14708 9764 15532
rect 8592 14680 9764 14708
rect 10004 15532 11176 15560
rect 10004 14708 11092 15532
rect 11156 14708 11176 15532
rect 10004 14680 11176 14708
rect 11416 15532 12588 15560
rect 11416 14708 12504 15532
rect 12568 14708 12588 15532
rect 11416 14680 12588 14708
rect 12828 15532 14000 15560
rect 12828 14708 13916 15532
rect 13980 14708 14000 15532
rect 12828 14680 14000 14708
rect 14240 15532 15412 15560
rect 14240 14708 15328 15532
rect 15392 14708 15412 15532
rect 14240 14680 15412 14708
rect 15652 15532 16824 15560
rect 15652 14708 16740 15532
rect 16804 14708 16824 15532
rect 15652 14680 16824 14708
rect 17064 15532 18236 15560
rect 17064 14708 18152 15532
rect 18216 14708 18236 15532
rect 17064 14680 18236 14708
rect 18476 15532 19648 15560
rect 18476 14708 19564 15532
rect 19628 14708 19648 15532
rect 18476 14680 19648 14708
rect 19888 15532 21060 15560
rect 19888 14708 20976 15532
rect 21040 14708 21060 15532
rect 19888 14680 21060 14708
rect 21300 15532 22472 15560
rect 21300 14708 22388 15532
rect 22452 14708 22472 15532
rect 21300 14680 22472 14708
rect 22712 15532 23884 15560
rect 22712 14708 23800 15532
rect 23864 14708 23884 15532
rect 22712 14680 23884 14708
rect -23884 14412 -22712 14440
rect -23884 13588 -22796 14412
rect -22732 13588 -22712 14412
rect -23884 13560 -22712 13588
rect -22472 14412 -21300 14440
rect -22472 13588 -21384 14412
rect -21320 13588 -21300 14412
rect -22472 13560 -21300 13588
rect -21060 14412 -19888 14440
rect -21060 13588 -19972 14412
rect -19908 13588 -19888 14412
rect -21060 13560 -19888 13588
rect -19648 14412 -18476 14440
rect -19648 13588 -18560 14412
rect -18496 13588 -18476 14412
rect -19648 13560 -18476 13588
rect -18236 14412 -17064 14440
rect -18236 13588 -17148 14412
rect -17084 13588 -17064 14412
rect -18236 13560 -17064 13588
rect -16824 14412 -15652 14440
rect -16824 13588 -15736 14412
rect -15672 13588 -15652 14412
rect -16824 13560 -15652 13588
rect -15412 14412 -14240 14440
rect -15412 13588 -14324 14412
rect -14260 13588 -14240 14412
rect -15412 13560 -14240 13588
rect -14000 14412 -12828 14440
rect -14000 13588 -12912 14412
rect -12848 13588 -12828 14412
rect -14000 13560 -12828 13588
rect -12588 14412 -11416 14440
rect -12588 13588 -11500 14412
rect -11436 13588 -11416 14412
rect -12588 13560 -11416 13588
rect -11176 14412 -10004 14440
rect -11176 13588 -10088 14412
rect -10024 13588 -10004 14412
rect -11176 13560 -10004 13588
rect -9764 14412 -8592 14440
rect -9764 13588 -8676 14412
rect -8612 13588 -8592 14412
rect -9764 13560 -8592 13588
rect -8352 14412 -7180 14440
rect -8352 13588 -7264 14412
rect -7200 13588 -7180 14412
rect -8352 13560 -7180 13588
rect -6940 14412 -5768 14440
rect -6940 13588 -5852 14412
rect -5788 13588 -5768 14412
rect -6940 13560 -5768 13588
rect -5528 14412 -4356 14440
rect -5528 13588 -4440 14412
rect -4376 13588 -4356 14412
rect -5528 13560 -4356 13588
rect -4116 14412 -2944 14440
rect -4116 13588 -3028 14412
rect -2964 13588 -2944 14412
rect -4116 13560 -2944 13588
rect -2704 14412 -1532 14440
rect -2704 13588 -1616 14412
rect -1552 13588 -1532 14412
rect -2704 13560 -1532 13588
rect -1292 14412 -120 14440
rect -1292 13588 -204 14412
rect -140 13588 -120 14412
rect -1292 13560 -120 13588
rect 120 14412 1292 14440
rect 120 13588 1208 14412
rect 1272 13588 1292 14412
rect 120 13560 1292 13588
rect 1532 14412 2704 14440
rect 1532 13588 2620 14412
rect 2684 13588 2704 14412
rect 1532 13560 2704 13588
rect 2944 14412 4116 14440
rect 2944 13588 4032 14412
rect 4096 13588 4116 14412
rect 2944 13560 4116 13588
rect 4356 14412 5528 14440
rect 4356 13588 5444 14412
rect 5508 13588 5528 14412
rect 4356 13560 5528 13588
rect 5768 14412 6940 14440
rect 5768 13588 6856 14412
rect 6920 13588 6940 14412
rect 5768 13560 6940 13588
rect 7180 14412 8352 14440
rect 7180 13588 8268 14412
rect 8332 13588 8352 14412
rect 7180 13560 8352 13588
rect 8592 14412 9764 14440
rect 8592 13588 9680 14412
rect 9744 13588 9764 14412
rect 8592 13560 9764 13588
rect 10004 14412 11176 14440
rect 10004 13588 11092 14412
rect 11156 13588 11176 14412
rect 10004 13560 11176 13588
rect 11416 14412 12588 14440
rect 11416 13588 12504 14412
rect 12568 13588 12588 14412
rect 11416 13560 12588 13588
rect 12828 14412 14000 14440
rect 12828 13588 13916 14412
rect 13980 13588 14000 14412
rect 12828 13560 14000 13588
rect 14240 14412 15412 14440
rect 14240 13588 15328 14412
rect 15392 13588 15412 14412
rect 14240 13560 15412 13588
rect 15652 14412 16824 14440
rect 15652 13588 16740 14412
rect 16804 13588 16824 14412
rect 15652 13560 16824 13588
rect 17064 14412 18236 14440
rect 17064 13588 18152 14412
rect 18216 13588 18236 14412
rect 17064 13560 18236 13588
rect 18476 14412 19648 14440
rect 18476 13588 19564 14412
rect 19628 13588 19648 14412
rect 18476 13560 19648 13588
rect 19888 14412 21060 14440
rect 19888 13588 20976 14412
rect 21040 13588 21060 14412
rect 19888 13560 21060 13588
rect 21300 14412 22472 14440
rect 21300 13588 22388 14412
rect 22452 13588 22472 14412
rect 21300 13560 22472 13588
rect 22712 14412 23884 14440
rect 22712 13588 23800 14412
rect 23864 13588 23884 14412
rect 22712 13560 23884 13588
rect -23884 13292 -22712 13320
rect -23884 12468 -22796 13292
rect -22732 12468 -22712 13292
rect -23884 12440 -22712 12468
rect -22472 13292 -21300 13320
rect -22472 12468 -21384 13292
rect -21320 12468 -21300 13292
rect -22472 12440 -21300 12468
rect -21060 13292 -19888 13320
rect -21060 12468 -19972 13292
rect -19908 12468 -19888 13292
rect -21060 12440 -19888 12468
rect -19648 13292 -18476 13320
rect -19648 12468 -18560 13292
rect -18496 12468 -18476 13292
rect -19648 12440 -18476 12468
rect -18236 13292 -17064 13320
rect -18236 12468 -17148 13292
rect -17084 12468 -17064 13292
rect -18236 12440 -17064 12468
rect -16824 13292 -15652 13320
rect -16824 12468 -15736 13292
rect -15672 12468 -15652 13292
rect -16824 12440 -15652 12468
rect -15412 13292 -14240 13320
rect -15412 12468 -14324 13292
rect -14260 12468 -14240 13292
rect -15412 12440 -14240 12468
rect -14000 13292 -12828 13320
rect -14000 12468 -12912 13292
rect -12848 12468 -12828 13292
rect -14000 12440 -12828 12468
rect -12588 13292 -11416 13320
rect -12588 12468 -11500 13292
rect -11436 12468 -11416 13292
rect -12588 12440 -11416 12468
rect -11176 13292 -10004 13320
rect -11176 12468 -10088 13292
rect -10024 12468 -10004 13292
rect -11176 12440 -10004 12468
rect -9764 13292 -8592 13320
rect -9764 12468 -8676 13292
rect -8612 12468 -8592 13292
rect -9764 12440 -8592 12468
rect -8352 13292 -7180 13320
rect -8352 12468 -7264 13292
rect -7200 12468 -7180 13292
rect -8352 12440 -7180 12468
rect -6940 13292 -5768 13320
rect -6940 12468 -5852 13292
rect -5788 12468 -5768 13292
rect -6940 12440 -5768 12468
rect -5528 13292 -4356 13320
rect -5528 12468 -4440 13292
rect -4376 12468 -4356 13292
rect -5528 12440 -4356 12468
rect -4116 13292 -2944 13320
rect -4116 12468 -3028 13292
rect -2964 12468 -2944 13292
rect -4116 12440 -2944 12468
rect -2704 13292 -1532 13320
rect -2704 12468 -1616 13292
rect -1552 12468 -1532 13292
rect -2704 12440 -1532 12468
rect -1292 13292 -120 13320
rect -1292 12468 -204 13292
rect -140 12468 -120 13292
rect -1292 12440 -120 12468
rect 120 13292 1292 13320
rect 120 12468 1208 13292
rect 1272 12468 1292 13292
rect 120 12440 1292 12468
rect 1532 13292 2704 13320
rect 1532 12468 2620 13292
rect 2684 12468 2704 13292
rect 1532 12440 2704 12468
rect 2944 13292 4116 13320
rect 2944 12468 4032 13292
rect 4096 12468 4116 13292
rect 2944 12440 4116 12468
rect 4356 13292 5528 13320
rect 4356 12468 5444 13292
rect 5508 12468 5528 13292
rect 4356 12440 5528 12468
rect 5768 13292 6940 13320
rect 5768 12468 6856 13292
rect 6920 12468 6940 13292
rect 5768 12440 6940 12468
rect 7180 13292 8352 13320
rect 7180 12468 8268 13292
rect 8332 12468 8352 13292
rect 7180 12440 8352 12468
rect 8592 13292 9764 13320
rect 8592 12468 9680 13292
rect 9744 12468 9764 13292
rect 8592 12440 9764 12468
rect 10004 13292 11176 13320
rect 10004 12468 11092 13292
rect 11156 12468 11176 13292
rect 10004 12440 11176 12468
rect 11416 13292 12588 13320
rect 11416 12468 12504 13292
rect 12568 12468 12588 13292
rect 11416 12440 12588 12468
rect 12828 13292 14000 13320
rect 12828 12468 13916 13292
rect 13980 12468 14000 13292
rect 12828 12440 14000 12468
rect 14240 13292 15412 13320
rect 14240 12468 15328 13292
rect 15392 12468 15412 13292
rect 14240 12440 15412 12468
rect 15652 13292 16824 13320
rect 15652 12468 16740 13292
rect 16804 12468 16824 13292
rect 15652 12440 16824 12468
rect 17064 13292 18236 13320
rect 17064 12468 18152 13292
rect 18216 12468 18236 13292
rect 17064 12440 18236 12468
rect 18476 13292 19648 13320
rect 18476 12468 19564 13292
rect 19628 12468 19648 13292
rect 18476 12440 19648 12468
rect 19888 13292 21060 13320
rect 19888 12468 20976 13292
rect 21040 12468 21060 13292
rect 19888 12440 21060 12468
rect 21300 13292 22472 13320
rect 21300 12468 22388 13292
rect 22452 12468 22472 13292
rect 21300 12440 22472 12468
rect 22712 13292 23884 13320
rect 22712 12468 23800 13292
rect 23864 12468 23884 13292
rect 22712 12440 23884 12468
rect -23884 12172 -22712 12200
rect -23884 11348 -22796 12172
rect -22732 11348 -22712 12172
rect -23884 11320 -22712 11348
rect -22472 12172 -21300 12200
rect -22472 11348 -21384 12172
rect -21320 11348 -21300 12172
rect -22472 11320 -21300 11348
rect -21060 12172 -19888 12200
rect -21060 11348 -19972 12172
rect -19908 11348 -19888 12172
rect -21060 11320 -19888 11348
rect -19648 12172 -18476 12200
rect -19648 11348 -18560 12172
rect -18496 11348 -18476 12172
rect -19648 11320 -18476 11348
rect -18236 12172 -17064 12200
rect -18236 11348 -17148 12172
rect -17084 11348 -17064 12172
rect -18236 11320 -17064 11348
rect -16824 12172 -15652 12200
rect -16824 11348 -15736 12172
rect -15672 11348 -15652 12172
rect -16824 11320 -15652 11348
rect -15412 12172 -14240 12200
rect -15412 11348 -14324 12172
rect -14260 11348 -14240 12172
rect -15412 11320 -14240 11348
rect -14000 12172 -12828 12200
rect -14000 11348 -12912 12172
rect -12848 11348 -12828 12172
rect -14000 11320 -12828 11348
rect -12588 12172 -11416 12200
rect -12588 11348 -11500 12172
rect -11436 11348 -11416 12172
rect -12588 11320 -11416 11348
rect -11176 12172 -10004 12200
rect -11176 11348 -10088 12172
rect -10024 11348 -10004 12172
rect -11176 11320 -10004 11348
rect -9764 12172 -8592 12200
rect -9764 11348 -8676 12172
rect -8612 11348 -8592 12172
rect -9764 11320 -8592 11348
rect -8352 12172 -7180 12200
rect -8352 11348 -7264 12172
rect -7200 11348 -7180 12172
rect -8352 11320 -7180 11348
rect -6940 12172 -5768 12200
rect -6940 11348 -5852 12172
rect -5788 11348 -5768 12172
rect -6940 11320 -5768 11348
rect -5528 12172 -4356 12200
rect -5528 11348 -4440 12172
rect -4376 11348 -4356 12172
rect -5528 11320 -4356 11348
rect -4116 12172 -2944 12200
rect -4116 11348 -3028 12172
rect -2964 11348 -2944 12172
rect -4116 11320 -2944 11348
rect -2704 12172 -1532 12200
rect -2704 11348 -1616 12172
rect -1552 11348 -1532 12172
rect -2704 11320 -1532 11348
rect -1292 12172 -120 12200
rect -1292 11348 -204 12172
rect -140 11348 -120 12172
rect -1292 11320 -120 11348
rect 120 12172 1292 12200
rect 120 11348 1208 12172
rect 1272 11348 1292 12172
rect 120 11320 1292 11348
rect 1532 12172 2704 12200
rect 1532 11348 2620 12172
rect 2684 11348 2704 12172
rect 1532 11320 2704 11348
rect 2944 12172 4116 12200
rect 2944 11348 4032 12172
rect 4096 11348 4116 12172
rect 2944 11320 4116 11348
rect 4356 12172 5528 12200
rect 4356 11348 5444 12172
rect 5508 11348 5528 12172
rect 4356 11320 5528 11348
rect 5768 12172 6940 12200
rect 5768 11348 6856 12172
rect 6920 11348 6940 12172
rect 5768 11320 6940 11348
rect 7180 12172 8352 12200
rect 7180 11348 8268 12172
rect 8332 11348 8352 12172
rect 7180 11320 8352 11348
rect 8592 12172 9764 12200
rect 8592 11348 9680 12172
rect 9744 11348 9764 12172
rect 8592 11320 9764 11348
rect 10004 12172 11176 12200
rect 10004 11348 11092 12172
rect 11156 11348 11176 12172
rect 10004 11320 11176 11348
rect 11416 12172 12588 12200
rect 11416 11348 12504 12172
rect 12568 11348 12588 12172
rect 11416 11320 12588 11348
rect 12828 12172 14000 12200
rect 12828 11348 13916 12172
rect 13980 11348 14000 12172
rect 12828 11320 14000 11348
rect 14240 12172 15412 12200
rect 14240 11348 15328 12172
rect 15392 11348 15412 12172
rect 14240 11320 15412 11348
rect 15652 12172 16824 12200
rect 15652 11348 16740 12172
rect 16804 11348 16824 12172
rect 15652 11320 16824 11348
rect 17064 12172 18236 12200
rect 17064 11348 18152 12172
rect 18216 11348 18236 12172
rect 17064 11320 18236 11348
rect 18476 12172 19648 12200
rect 18476 11348 19564 12172
rect 19628 11348 19648 12172
rect 18476 11320 19648 11348
rect 19888 12172 21060 12200
rect 19888 11348 20976 12172
rect 21040 11348 21060 12172
rect 19888 11320 21060 11348
rect 21300 12172 22472 12200
rect 21300 11348 22388 12172
rect 22452 11348 22472 12172
rect 21300 11320 22472 11348
rect 22712 12172 23884 12200
rect 22712 11348 23800 12172
rect 23864 11348 23884 12172
rect 22712 11320 23884 11348
rect -23884 11052 -22712 11080
rect -23884 10228 -22796 11052
rect -22732 10228 -22712 11052
rect -23884 10200 -22712 10228
rect -22472 11052 -21300 11080
rect -22472 10228 -21384 11052
rect -21320 10228 -21300 11052
rect -22472 10200 -21300 10228
rect -21060 11052 -19888 11080
rect -21060 10228 -19972 11052
rect -19908 10228 -19888 11052
rect -21060 10200 -19888 10228
rect -19648 11052 -18476 11080
rect -19648 10228 -18560 11052
rect -18496 10228 -18476 11052
rect -19648 10200 -18476 10228
rect -18236 11052 -17064 11080
rect -18236 10228 -17148 11052
rect -17084 10228 -17064 11052
rect -18236 10200 -17064 10228
rect -16824 11052 -15652 11080
rect -16824 10228 -15736 11052
rect -15672 10228 -15652 11052
rect -16824 10200 -15652 10228
rect -15412 11052 -14240 11080
rect -15412 10228 -14324 11052
rect -14260 10228 -14240 11052
rect -15412 10200 -14240 10228
rect -14000 11052 -12828 11080
rect -14000 10228 -12912 11052
rect -12848 10228 -12828 11052
rect -14000 10200 -12828 10228
rect -12588 11052 -11416 11080
rect -12588 10228 -11500 11052
rect -11436 10228 -11416 11052
rect -12588 10200 -11416 10228
rect -11176 11052 -10004 11080
rect -11176 10228 -10088 11052
rect -10024 10228 -10004 11052
rect -11176 10200 -10004 10228
rect -9764 11052 -8592 11080
rect -9764 10228 -8676 11052
rect -8612 10228 -8592 11052
rect -9764 10200 -8592 10228
rect -8352 11052 -7180 11080
rect -8352 10228 -7264 11052
rect -7200 10228 -7180 11052
rect -8352 10200 -7180 10228
rect -6940 11052 -5768 11080
rect -6940 10228 -5852 11052
rect -5788 10228 -5768 11052
rect -6940 10200 -5768 10228
rect -5528 11052 -4356 11080
rect -5528 10228 -4440 11052
rect -4376 10228 -4356 11052
rect -5528 10200 -4356 10228
rect -4116 11052 -2944 11080
rect -4116 10228 -3028 11052
rect -2964 10228 -2944 11052
rect -4116 10200 -2944 10228
rect -2704 11052 -1532 11080
rect -2704 10228 -1616 11052
rect -1552 10228 -1532 11052
rect -2704 10200 -1532 10228
rect -1292 11052 -120 11080
rect -1292 10228 -204 11052
rect -140 10228 -120 11052
rect -1292 10200 -120 10228
rect 120 11052 1292 11080
rect 120 10228 1208 11052
rect 1272 10228 1292 11052
rect 120 10200 1292 10228
rect 1532 11052 2704 11080
rect 1532 10228 2620 11052
rect 2684 10228 2704 11052
rect 1532 10200 2704 10228
rect 2944 11052 4116 11080
rect 2944 10228 4032 11052
rect 4096 10228 4116 11052
rect 2944 10200 4116 10228
rect 4356 11052 5528 11080
rect 4356 10228 5444 11052
rect 5508 10228 5528 11052
rect 4356 10200 5528 10228
rect 5768 11052 6940 11080
rect 5768 10228 6856 11052
rect 6920 10228 6940 11052
rect 5768 10200 6940 10228
rect 7180 11052 8352 11080
rect 7180 10228 8268 11052
rect 8332 10228 8352 11052
rect 7180 10200 8352 10228
rect 8592 11052 9764 11080
rect 8592 10228 9680 11052
rect 9744 10228 9764 11052
rect 8592 10200 9764 10228
rect 10004 11052 11176 11080
rect 10004 10228 11092 11052
rect 11156 10228 11176 11052
rect 10004 10200 11176 10228
rect 11416 11052 12588 11080
rect 11416 10228 12504 11052
rect 12568 10228 12588 11052
rect 11416 10200 12588 10228
rect 12828 11052 14000 11080
rect 12828 10228 13916 11052
rect 13980 10228 14000 11052
rect 12828 10200 14000 10228
rect 14240 11052 15412 11080
rect 14240 10228 15328 11052
rect 15392 10228 15412 11052
rect 14240 10200 15412 10228
rect 15652 11052 16824 11080
rect 15652 10228 16740 11052
rect 16804 10228 16824 11052
rect 15652 10200 16824 10228
rect 17064 11052 18236 11080
rect 17064 10228 18152 11052
rect 18216 10228 18236 11052
rect 17064 10200 18236 10228
rect 18476 11052 19648 11080
rect 18476 10228 19564 11052
rect 19628 10228 19648 11052
rect 18476 10200 19648 10228
rect 19888 11052 21060 11080
rect 19888 10228 20976 11052
rect 21040 10228 21060 11052
rect 19888 10200 21060 10228
rect 21300 11052 22472 11080
rect 21300 10228 22388 11052
rect 22452 10228 22472 11052
rect 21300 10200 22472 10228
rect 22712 11052 23884 11080
rect 22712 10228 23800 11052
rect 23864 10228 23884 11052
rect 22712 10200 23884 10228
rect -23884 9932 -22712 9960
rect -23884 9108 -22796 9932
rect -22732 9108 -22712 9932
rect -23884 9080 -22712 9108
rect -22472 9932 -21300 9960
rect -22472 9108 -21384 9932
rect -21320 9108 -21300 9932
rect -22472 9080 -21300 9108
rect -21060 9932 -19888 9960
rect -21060 9108 -19972 9932
rect -19908 9108 -19888 9932
rect -21060 9080 -19888 9108
rect -19648 9932 -18476 9960
rect -19648 9108 -18560 9932
rect -18496 9108 -18476 9932
rect -19648 9080 -18476 9108
rect -18236 9932 -17064 9960
rect -18236 9108 -17148 9932
rect -17084 9108 -17064 9932
rect -18236 9080 -17064 9108
rect -16824 9932 -15652 9960
rect -16824 9108 -15736 9932
rect -15672 9108 -15652 9932
rect -16824 9080 -15652 9108
rect -15412 9932 -14240 9960
rect -15412 9108 -14324 9932
rect -14260 9108 -14240 9932
rect -15412 9080 -14240 9108
rect -14000 9932 -12828 9960
rect -14000 9108 -12912 9932
rect -12848 9108 -12828 9932
rect -14000 9080 -12828 9108
rect -12588 9932 -11416 9960
rect -12588 9108 -11500 9932
rect -11436 9108 -11416 9932
rect -12588 9080 -11416 9108
rect -11176 9932 -10004 9960
rect -11176 9108 -10088 9932
rect -10024 9108 -10004 9932
rect -11176 9080 -10004 9108
rect -9764 9932 -8592 9960
rect -9764 9108 -8676 9932
rect -8612 9108 -8592 9932
rect -9764 9080 -8592 9108
rect -8352 9932 -7180 9960
rect -8352 9108 -7264 9932
rect -7200 9108 -7180 9932
rect -8352 9080 -7180 9108
rect -6940 9932 -5768 9960
rect -6940 9108 -5852 9932
rect -5788 9108 -5768 9932
rect -6940 9080 -5768 9108
rect -5528 9932 -4356 9960
rect -5528 9108 -4440 9932
rect -4376 9108 -4356 9932
rect -5528 9080 -4356 9108
rect -4116 9932 -2944 9960
rect -4116 9108 -3028 9932
rect -2964 9108 -2944 9932
rect -4116 9080 -2944 9108
rect -2704 9932 -1532 9960
rect -2704 9108 -1616 9932
rect -1552 9108 -1532 9932
rect -2704 9080 -1532 9108
rect -1292 9932 -120 9960
rect -1292 9108 -204 9932
rect -140 9108 -120 9932
rect -1292 9080 -120 9108
rect 120 9932 1292 9960
rect 120 9108 1208 9932
rect 1272 9108 1292 9932
rect 120 9080 1292 9108
rect 1532 9932 2704 9960
rect 1532 9108 2620 9932
rect 2684 9108 2704 9932
rect 1532 9080 2704 9108
rect 2944 9932 4116 9960
rect 2944 9108 4032 9932
rect 4096 9108 4116 9932
rect 2944 9080 4116 9108
rect 4356 9932 5528 9960
rect 4356 9108 5444 9932
rect 5508 9108 5528 9932
rect 4356 9080 5528 9108
rect 5768 9932 6940 9960
rect 5768 9108 6856 9932
rect 6920 9108 6940 9932
rect 5768 9080 6940 9108
rect 7180 9932 8352 9960
rect 7180 9108 8268 9932
rect 8332 9108 8352 9932
rect 7180 9080 8352 9108
rect 8592 9932 9764 9960
rect 8592 9108 9680 9932
rect 9744 9108 9764 9932
rect 8592 9080 9764 9108
rect 10004 9932 11176 9960
rect 10004 9108 11092 9932
rect 11156 9108 11176 9932
rect 10004 9080 11176 9108
rect 11416 9932 12588 9960
rect 11416 9108 12504 9932
rect 12568 9108 12588 9932
rect 11416 9080 12588 9108
rect 12828 9932 14000 9960
rect 12828 9108 13916 9932
rect 13980 9108 14000 9932
rect 12828 9080 14000 9108
rect 14240 9932 15412 9960
rect 14240 9108 15328 9932
rect 15392 9108 15412 9932
rect 14240 9080 15412 9108
rect 15652 9932 16824 9960
rect 15652 9108 16740 9932
rect 16804 9108 16824 9932
rect 15652 9080 16824 9108
rect 17064 9932 18236 9960
rect 17064 9108 18152 9932
rect 18216 9108 18236 9932
rect 17064 9080 18236 9108
rect 18476 9932 19648 9960
rect 18476 9108 19564 9932
rect 19628 9108 19648 9932
rect 18476 9080 19648 9108
rect 19888 9932 21060 9960
rect 19888 9108 20976 9932
rect 21040 9108 21060 9932
rect 19888 9080 21060 9108
rect 21300 9932 22472 9960
rect 21300 9108 22388 9932
rect 22452 9108 22472 9932
rect 21300 9080 22472 9108
rect 22712 9932 23884 9960
rect 22712 9108 23800 9932
rect 23864 9108 23884 9932
rect 22712 9080 23884 9108
rect -23884 8812 -22712 8840
rect -23884 7988 -22796 8812
rect -22732 7988 -22712 8812
rect -23884 7960 -22712 7988
rect -22472 8812 -21300 8840
rect -22472 7988 -21384 8812
rect -21320 7988 -21300 8812
rect -22472 7960 -21300 7988
rect -21060 8812 -19888 8840
rect -21060 7988 -19972 8812
rect -19908 7988 -19888 8812
rect -21060 7960 -19888 7988
rect -19648 8812 -18476 8840
rect -19648 7988 -18560 8812
rect -18496 7988 -18476 8812
rect -19648 7960 -18476 7988
rect -18236 8812 -17064 8840
rect -18236 7988 -17148 8812
rect -17084 7988 -17064 8812
rect -18236 7960 -17064 7988
rect -16824 8812 -15652 8840
rect -16824 7988 -15736 8812
rect -15672 7988 -15652 8812
rect -16824 7960 -15652 7988
rect -15412 8812 -14240 8840
rect -15412 7988 -14324 8812
rect -14260 7988 -14240 8812
rect -15412 7960 -14240 7988
rect -14000 8812 -12828 8840
rect -14000 7988 -12912 8812
rect -12848 7988 -12828 8812
rect -14000 7960 -12828 7988
rect -12588 8812 -11416 8840
rect -12588 7988 -11500 8812
rect -11436 7988 -11416 8812
rect -12588 7960 -11416 7988
rect -11176 8812 -10004 8840
rect -11176 7988 -10088 8812
rect -10024 7988 -10004 8812
rect -11176 7960 -10004 7988
rect -9764 8812 -8592 8840
rect -9764 7988 -8676 8812
rect -8612 7988 -8592 8812
rect -9764 7960 -8592 7988
rect -8352 8812 -7180 8840
rect -8352 7988 -7264 8812
rect -7200 7988 -7180 8812
rect -8352 7960 -7180 7988
rect -6940 8812 -5768 8840
rect -6940 7988 -5852 8812
rect -5788 7988 -5768 8812
rect -6940 7960 -5768 7988
rect -5528 8812 -4356 8840
rect -5528 7988 -4440 8812
rect -4376 7988 -4356 8812
rect -5528 7960 -4356 7988
rect -4116 8812 -2944 8840
rect -4116 7988 -3028 8812
rect -2964 7988 -2944 8812
rect -4116 7960 -2944 7988
rect -2704 8812 -1532 8840
rect -2704 7988 -1616 8812
rect -1552 7988 -1532 8812
rect -2704 7960 -1532 7988
rect -1292 8812 -120 8840
rect -1292 7988 -204 8812
rect -140 7988 -120 8812
rect -1292 7960 -120 7988
rect 120 8812 1292 8840
rect 120 7988 1208 8812
rect 1272 7988 1292 8812
rect 120 7960 1292 7988
rect 1532 8812 2704 8840
rect 1532 7988 2620 8812
rect 2684 7988 2704 8812
rect 1532 7960 2704 7988
rect 2944 8812 4116 8840
rect 2944 7988 4032 8812
rect 4096 7988 4116 8812
rect 2944 7960 4116 7988
rect 4356 8812 5528 8840
rect 4356 7988 5444 8812
rect 5508 7988 5528 8812
rect 4356 7960 5528 7988
rect 5768 8812 6940 8840
rect 5768 7988 6856 8812
rect 6920 7988 6940 8812
rect 5768 7960 6940 7988
rect 7180 8812 8352 8840
rect 7180 7988 8268 8812
rect 8332 7988 8352 8812
rect 7180 7960 8352 7988
rect 8592 8812 9764 8840
rect 8592 7988 9680 8812
rect 9744 7988 9764 8812
rect 8592 7960 9764 7988
rect 10004 8812 11176 8840
rect 10004 7988 11092 8812
rect 11156 7988 11176 8812
rect 10004 7960 11176 7988
rect 11416 8812 12588 8840
rect 11416 7988 12504 8812
rect 12568 7988 12588 8812
rect 11416 7960 12588 7988
rect 12828 8812 14000 8840
rect 12828 7988 13916 8812
rect 13980 7988 14000 8812
rect 12828 7960 14000 7988
rect 14240 8812 15412 8840
rect 14240 7988 15328 8812
rect 15392 7988 15412 8812
rect 14240 7960 15412 7988
rect 15652 8812 16824 8840
rect 15652 7988 16740 8812
rect 16804 7988 16824 8812
rect 15652 7960 16824 7988
rect 17064 8812 18236 8840
rect 17064 7988 18152 8812
rect 18216 7988 18236 8812
rect 17064 7960 18236 7988
rect 18476 8812 19648 8840
rect 18476 7988 19564 8812
rect 19628 7988 19648 8812
rect 18476 7960 19648 7988
rect 19888 8812 21060 8840
rect 19888 7988 20976 8812
rect 21040 7988 21060 8812
rect 19888 7960 21060 7988
rect 21300 8812 22472 8840
rect 21300 7988 22388 8812
rect 22452 7988 22472 8812
rect 21300 7960 22472 7988
rect 22712 8812 23884 8840
rect 22712 7988 23800 8812
rect 23864 7988 23884 8812
rect 22712 7960 23884 7988
rect -23884 7692 -22712 7720
rect -23884 6868 -22796 7692
rect -22732 6868 -22712 7692
rect -23884 6840 -22712 6868
rect -22472 7692 -21300 7720
rect -22472 6868 -21384 7692
rect -21320 6868 -21300 7692
rect -22472 6840 -21300 6868
rect -21060 7692 -19888 7720
rect -21060 6868 -19972 7692
rect -19908 6868 -19888 7692
rect -21060 6840 -19888 6868
rect -19648 7692 -18476 7720
rect -19648 6868 -18560 7692
rect -18496 6868 -18476 7692
rect -19648 6840 -18476 6868
rect -18236 7692 -17064 7720
rect -18236 6868 -17148 7692
rect -17084 6868 -17064 7692
rect -18236 6840 -17064 6868
rect -16824 7692 -15652 7720
rect -16824 6868 -15736 7692
rect -15672 6868 -15652 7692
rect -16824 6840 -15652 6868
rect -15412 7692 -14240 7720
rect -15412 6868 -14324 7692
rect -14260 6868 -14240 7692
rect -15412 6840 -14240 6868
rect -14000 7692 -12828 7720
rect -14000 6868 -12912 7692
rect -12848 6868 -12828 7692
rect -14000 6840 -12828 6868
rect -12588 7692 -11416 7720
rect -12588 6868 -11500 7692
rect -11436 6868 -11416 7692
rect -12588 6840 -11416 6868
rect -11176 7692 -10004 7720
rect -11176 6868 -10088 7692
rect -10024 6868 -10004 7692
rect -11176 6840 -10004 6868
rect -9764 7692 -8592 7720
rect -9764 6868 -8676 7692
rect -8612 6868 -8592 7692
rect -9764 6840 -8592 6868
rect -8352 7692 -7180 7720
rect -8352 6868 -7264 7692
rect -7200 6868 -7180 7692
rect -8352 6840 -7180 6868
rect -6940 7692 -5768 7720
rect -6940 6868 -5852 7692
rect -5788 6868 -5768 7692
rect -6940 6840 -5768 6868
rect -5528 7692 -4356 7720
rect -5528 6868 -4440 7692
rect -4376 6868 -4356 7692
rect -5528 6840 -4356 6868
rect -4116 7692 -2944 7720
rect -4116 6868 -3028 7692
rect -2964 6868 -2944 7692
rect -4116 6840 -2944 6868
rect -2704 7692 -1532 7720
rect -2704 6868 -1616 7692
rect -1552 6868 -1532 7692
rect -2704 6840 -1532 6868
rect -1292 7692 -120 7720
rect -1292 6868 -204 7692
rect -140 6868 -120 7692
rect -1292 6840 -120 6868
rect 120 7692 1292 7720
rect 120 6868 1208 7692
rect 1272 6868 1292 7692
rect 120 6840 1292 6868
rect 1532 7692 2704 7720
rect 1532 6868 2620 7692
rect 2684 6868 2704 7692
rect 1532 6840 2704 6868
rect 2944 7692 4116 7720
rect 2944 6868 4032 7692
rect 4096 6868 4116 7692
rect 2944 6840 4116 6868
rect 4356 7692 5528 7720
rect 4356 6868 5444 7692
rect 5508 6868 5528 7692
rect 4356 6840 5528 6868
rect 5768 7692 6940 7720
rect 5768 6868 6856 7692
rect 6920 6868 6940 7692
rect 5768 6840 6940 6868
rect 7180 7692 8352 7720
rect 7180 6868 8268 7692
rect 8332 6868 8352 7692
rect 7180 6840 8352 6868
rect 8592 7692 9764 7720
rect 8592 6868 9680 7692
rect 9744 6868 9764 7692
rect 8592 6840 9764 6868
rect 10004 7692 11176 7720
rect 10004 6868 11092 7692
rect 11156 6868 11176 7692
rect 10004 6840 11176 6868
rect 11416 7692 12588 7720
rect 11416 6868 12504 7692
rect 12568 6868 12588 7692
rect 11416 6840 12588 6868
rect 12828 7692 14000 7720
rect 12828 6868 13916 7692
rect 13980 6868 14000 7692
rect 12828 6840 14000 6868
rect 14240 7692 15412 7720
rect 14240 6868 15328 7692
rect 15392 6868 15412 7692
rect 14240 6840 15412 6868
rect 15652 7692 16824 7720
rect 15652 6868 16740 7692
rect 16804 6868 16824 7692
rect 15652 6840 16824 6868
rect 17064 7692 18236 7720
rect 17064 6868 18152 7692
rect 18216 6868 18236 7692
rect 17064 6840 18236 6868
rect 18476 7692 19648 7720
rect 18476 6868 19564 7692
rect 19628 6868 19648 7692
rect 18476 6840 19648 6868
rect 19888 7692 21060 7720
rect 19888 6868 20976 7692
rect 21040 6868 21060 7692
rect 19888 6840 21060 6868
rect 21300 7692 22472 7720
rect 21300 6868 22388 7692
rect 22452 6868 22472 7692
rect 21300 6840 22472 6868
rect 22712 7692 23884 7720
rect 22712 6868 23800 7692
rect 23864 6868 23884 7692
rect 22712 6840 23884 6868
rect -23884 6572 -22712 6600
rect -23884 5748 -22796 6572
rect -22732 5748 -22712 6572
rect -23884 5720 -22712 5748
rect -22472 6572 -21300 6600
rect -22472 5748 -21384 6572
rect -21320 5748 -21300 6572
rect -22472 5720 -21300 5748
rect -21060 6572 -19888 6600
rect -21060 5748 -19972 6572
rect -19908 5748 -19888 6572
rect -21060 5720 -19888 5748
rect -19648 6572 -18476 6600
rect -19648 5748 -18560 6572
rect -18496 5748 -18476 6572
rect -19648 5720 -18476 5748
rect -18236 6572 -17064 6600
rect -18236 5748 -17148 6572
rect -17084 5748 -17064 6572
rect -18236 5720 -17064 5748
rect -16824 6572 -15652 6600
rect -16824 5748 -15736 6572
rect -15672 5748 -15652 6572
rect -16824 5720 -15652 5748
rect -15412 6572 -14240 6600
rect -15412 5748 -14324 6572
rect -14260 5748 -14240 6572
rect -15412 5720 -14240 5748
rect -14000 6572 -12828 6600
rect -14000 5748 -12912 6572
rect -12848 5748 -12828 6572
rect -14000 5720 -12828 5748
rect -12588 6572 -11416 6600
rect -12588 5748 -11500 6572
rect -11436 5748 -11416 6572
rect -12588 5720 -11416 5748
rect -11176 6572 -10004 6600
rect -11176 5748 -10088 6572
rect -10024 5748 -10004 6572
rect -11176 5720 -10004 5748
rect -9764 6572 -8592 6600
rect -9764 5748 -8676 6572
rect -8612 5748 -8592 6572
rect -9764 5720 -8592 5748
rect -8352 6572 -7180 6600
rect -8352 5748 -7264 6572
rect -7200 5748 -7180 6572
rect -8352 5720 -7180 5748
rect -6940 6572 -5768 6600
rect -6940 5748 -5852 6572
rect -5788 5748 -5768 6572
rect -6940 5720 -5768 5748
rect -5528 6572 -4356 6600
rect -5528 5748 -4440 6572
rect -4376 5748 -4356 6572
rect -5528 5720 -4356 5748
rect -4116 6572 -2944 6600
rect -4116 5748 -3028 6572
rect -2964 5748 -2944 6572
rect -4116 5720 -2944 5748
rect -2704 6572 -1532 6600
rect -2704 5748 -1616 6572
rect -1552 5748 -1532 6572
rect -2704 5720 -1532 5748
rect -1292 6572 -120 6600
rect -1292 5748 -204 6572
rect -140 5748 -120 6572
rect -1292 5720 -120 5748
rect 120 6572 1292 6600
rect 120 5748 1208 6572
rect 1272 5748 1292 6572
rect 120 5720 1292 5748
rect 1532 6572 2704 6600
rect 1532 5748 2620 6572
rect 2684 5748 2704 6572
rect 1532 5720 2704 5748
rect 2944 6572 4116 6600
rect 2944 5748 4032 6572
rect 4096 5748 4116 6572
rect 2944 5720 4116 5748
rect 4356 6572 5528 6600
rect 4356 5748 5444 6572
rect 5508 5748 5528 6572
rect 4356 5720 5528 5748
rect 5768 6572 6940 6600
rect 5768 5748 6856 6572
rect 6920 5748 6940 6572
rect 5768 5720 6940 5748
rect 7180 6572 8352 6600
rect 7180 5748 8268 6572
rect 8332 5748 8352 6572
rect 7180 5720 8352 5748
rect 8592 6572 9764 6600
rect 8592 5748 9680 6572
rect 9744 5748 9764 6572
rect 8592 5720 9764 5748
rect 10004 6572 11176 6600
rect 10004 5748 11092 6572
rect 11156 5748 11176 6572
rect 10004 5720 11176 5748
rect 11416 6572 12588 6600
rect 11416 5748 12504 6572
rect 12568 5748 12588 6572
rect 11416 5720 12588 5748
rect 12828 6572 14000 6600
rect 12828 5748 13916 6572
rect 13980 5748 14000 6572
rect 12828 5720 14000 5748
rect 14240 6572 15412 6600
rect 14240 5748 15328 6572
rect 15392 5748 15412 6572
rect 14240 5720 15412 5748
rect 15652 6572 16824 6600
rect 15652 5748 16740 6572
rect 16804 5748 16824 6572
rect 15652 5720 16824 5748
rect 17064 6572 18236 6600
rect 17064 5748 18152 6572
rect 18216 5748 18236 6572
rect 17064 5720 18236 5748
rect 18476 6572 19648 6600
rect 18476 5748 19564 6572
rect 19628 5748 19648 6572
rect 18476 5720 19648 5748
rect 19888 6572 21060 6600
rect 19888 5748 20976 6572
rect 21040 5748 21060 6572
rect 19888 5720 21060 5748
rect 21300 6572 22472 6600
rect 21300 5748 22388 6572
rect 22452 5748 22472 6572
rect 21300 5720 22472 5748
rect 22712 6572 23884 6600
rect 22712 5748 23800 6572
rect 23864 5748 23884 6572
rect 22712 5720 23884 5748
rect -23884 5452 -22712 5480
rect -23884 4628 -22796 5452
rect -22732 4628 -22712 5452
rect -23884 4600 -22712 4628
rect -22472 5452 -21300 5480
rect -22472 4628 -21384 5452
rect -21320 4628 -21300 5452
rect -22472 4600 -21300 4628
rect -21060 5452 -19888 5480
rect -21060 4628 -19972 5452
rect -19908 4628 -19888 5452
rect -21060 4600 -19888 4628
rect -19648 5452 -18476 5480
rect -19648 4628 -18560 5452
rect -18496 4628 -18476 5452
rect -19648 4600 -18476 4628
rect -18236 5452 -17064 5480
rect -18236 4628 -17148 5452
rect -17084 4628 -17064 5452
rect -18236 4600 -17064 4628
rect -16824 5452 -15652 5480
rect -16824 4628 -15736 5452
rect -15672 4628 -15652 5452
rect -16824 4600 -15652 4628
rect -15412 5452 -14240 5480
rect -15412 4628 -14324 5452
rect -14260 4628 -14240 5452
rect -15412 4600 -14240 4628
rect -14000 5452 -12828 5480
rect -14000 4628 -12912 5452
rect -12848 4628 -12828 5452
rect -14000 4600 -12828 4628
rect -12588 5452 -11416 5480
rect -12588 4628 -11500 5452
rect -11436 4628 -11416 5452
rect -12588 4600 -11416 4628
rect -11176 5452 -10004 5480
rect -11176 4628 -10088 5452
rect -10024 4628 -10004 5452
rect -11176 4600 -10004 4628
rect -9764 5452 -8592 5480
rect -9764 4628 -8676 5452
rect -8612 4628 -8592 5452
rect -9764 4600 -8592 4628
rect -8352 5452 -7180 5480
rect -8352 4628 -7264 5452
rect -7200 4628 -7180 5452
rect -8352 4600 -7180 4628
rect -6940 5452 -5768 5480
rect -6940 4628 -5852 5452
rect -5788 4628 -5768 5452
rect -6940 4600 -5768 4628
rect -5528 5452 -4356 5480
rect -5528 4628 -4440 5452
rect -4376 4628 -4356 5452
rect -5528 4600 -4356 4628
rect -4116 5452 -2944 5480
rect -4116 4628 -3028 5452
rect -2964 4628 -2944 5452
rect -4116 4600 -2944 4628
rect -2704 5452 -1532 5480
rect -2704 4628 -1616 5452
rect -1552 4628 -1532 5452
rect -2704 4600 -1532 4628
rect -1292 5452 -120 5480
rect -1292 4628 -204 5452
rect -140 4628 -120 5452
rect -1292 4600 -120 4628
rect 120 5452 1292 5480
rect 120 4628 1208 5452
rect 1272 4628 1292 5452
rect 120 4600 1292 4628
rect 1532 5452 2704 5480
rect 1532 4628 2620 5452
rect 2684 4628 2704 5452
rect 1532 4600 2704 4628
rect 2944 5452 4116 5480
rect 2944 4628 4032 5452
rect 4096 4628 4116 5452
rect 2944 4600 4116 4628
rect 4356 5452 5528 5480
rect 4356 4628 5444 5452
rect 5508 4628 5528 5452
rect 4356 4600 5528 4628
rect 5768 5452 6940 5480
rect 5768 4628 6856 5452
rect 6920 4628 6940 5452
rect 5768 4600 6940 4628
rect 7180 5452 8352 5480
rect 7180 4628 8268 5452
rect 8332 4628 8352 5452
rect 7180 4600 8352 4628
rect 8592 5452 9764 5480
rect 8592 4628 9680 5452
rect 9744 4628 9764 5452
rect 8592 4600 9764 4628
rect 10004 5452 11176 5480
rect 10004 4628 11092 5452
rect 11156 4628 11176 5452
rect 10004 4600 11176 4628
rect 11416 5452 12588 5480
rect 11416 4628 12504 5452
rect 12568 4628 12588 5452
rect 11416 4600 12588 4628
rect 12828 5452 14000 5480
rect 12828 4628 13916 5452
rect 13980 4628 14000 5452
rect 12828 4600 14000 4628
rect 14240 5452 15412 5480
rect 14240 4628 15328 5452
rect 15392 4628 15412 5452
rect 14240 4600 15412 4628
rect 15652 5452 16824 5480
rect 15652 4628 16740 5452
rect 16804 4628 16824 5452
rect 15652 4600 16824 4628
rect 17064 5452 18236 5480
rect 17064 4628 18152 5452
rect 18216 4628 18236 5452
rect 17064 4600 18236 4628
rect 18476 5452 19648 5480
rect 18476 4628 19564 5452
rect 19628 4628 19648 5452
rect 18476 4600 19648 4628
rect 19888 5452 21060 5480
rect 19888 4628 20976 5452
rect 21040 4628 21060 5452
rect 19888 4600 21060 4628
rect 21300 5452 22472 5480
rect 21300 4628 22388 5452
rect 22452 4628 22472 5452
rect 21300 4600 22472 4628
rect 22712 5452 23884 5480
rect 22712 4628 23800 5452
rect 23864 4628 23884 5452
rect 22712 4600 23884 4628
rect -23884 4332 -22712 4360
rect -23884 3508 -22796 4332
rect -22732 3508 -22712 4332
rect -23884 3480 -22712 3508
rect -22472 4332 -21300 4360
rect -22472 3508 -21384 4332
rect -21320 3508 -21300 4332
rect -22472 3480 -21300 3508
rect -21060 4332 -19888 4360
rect -21060 3508 -19972 4332
rect -19908 3508 -19888 4332
rect -21060 3480 -19888 3508
rect -19648 4332 -18476 4360
rect -19648 3508 -18560 4332
rect -18496 3508 -18476 4332
rect -19648 3480 -18476 3508
rect -18236 4332 -17064 4360
rect -18236 3508 -17148 4332
rect -17084 3508 -17064 4332
rect -18236 3480 -17064 3508
rect -16824 4332 -15652 4360
rect -16824 3508 -15736 4332
rect -15672 3508 -15652 4332
rect -16824 3480 -15652 3508
rect -15412 4332 -14240 4360
rect -15412 3508 -14324 4332
rect -14260 3508 -14240 4332
rect -15412 3480 -14240 3508
rect -14000 4332 -12828 4360
rect -14000 3508 -12912 4332
rect -12848 3508 -12828 4332
rect -14000 3480 -12828 3508
rect -12588 4332 -11416 4360
rect -12588 3508 -11500 4332
rect -11436 3508 -11416 4332
rect -12588 3480 -11416 3508
rect -11176 4332 -10004 4360
rect -11176 3508 -10088 4332
rect -10024 3508 -10004 4332
rect -11176 3480 -10004 3508
rect -9764 4332 -8592 4360
rect -9764 3508 -8676 4332
rect -8612 3508 -8592 4332
rect -9764 3480 -8592 3508
rect -8352 4332 -7180 4360
rect -8352 3508 -7264 4332
rect -7200 3508 -7180 4332
rect -8352 3480 -7180 3508
rect -6940 4332 -5768 4360
rect -6940 3508 -5852 4332
rect -5788 3508 -5768 4332
rect -6940 3480 -5768 3508
rect -5528 4332 -4356 4360
rect -5528 3508 -4440 4332
rect -4376 3508 -4356 4332
rect -5528 3480 -4356 3508
rect -4116 4332 -2944 4360
rect -4116 3508 -3028 4332
rect -2964 3508 -2944 4332
rect -4116 3480 -2944 3508
rect -2704 4332 -1532 4360
rect -2704 3508 -1616 4332
rect -1552 3508 -1532 4332
rect -2704 3480 -1532 3508
rect -1292 4332 -120 4360
rect -1292 3508 -204 4332
rect -140 3508 -120 4332
rect -1292 3480 -120 3508
rect 120 4332 1292 4360
rect 120 3508 1208 4332
rect 1272 3508 1292 4332
rect 120 3480 1292 3508
rect 1532 4332 2704 4360
rect 1532 3508 2620 4332
rect 2684 3508 2704 4332
rect 1532 3480 2704 3508
rect 2944 4332 4116 4360
rect 2944 3508 4032 4332
rect 4096 3508 4116 4332
rect 2944 3480 4116 3508
rect 4356 4332 5528 4360
rect 4356 3508 5444 4332
rect 5508 3508 5528 4332
rect 4356 3480 5528 3508
rect 5768 4332 6940 4360
rect 5768 3508 6856 4332
rect 6920 3508 6940 4332
rect 5768 3480 6940 3508
rect 7180 4332 8352 4360
rect 7180 3508 8268 4332
rect 8332 3508 8352 4332
rect 7180 3480 8352 3508
rect 8592 4332 9764 4360
rect 8592 3508 9680 4332
rect 9744 3508 9764 4332
rect 8592 3480 9764 3508
rect 10004 4332 11176 4360
rect 10004 3508 11092 4332
rect 11156 3508 11176 4332
rect 10004 3480 11176 3508
rect 11416 4332 12588 4360
rect 11416 3508 12504 4332
rect 12568 3508 12588 4332
rect 11416 3480 12588 3508
rect 12828 4332 14000 4360
rect 12828 3508 13916 4332
rect 13980 3508 14000 4332
rect 12828 3480 14000 3508
rect 14240 4332 15412 4360
rect 14240 3508 15328 4332
rect 15392 3508 15412 4332
rect 14240 3480 15412 3508
rect 15652 4332 16824 4360
rect 15652 3508 16740 4332
rect 16804 3508 16824 4332
rect 15652 3480 16824 3508
rect 17064 4332 18236 4360
rect 17064 3508 18152 4332
rect 18216 3508 18236 4332
rect 17064 3480 18236 3508
rect 18476 4332 19648 4360
rect 18476 3508 19564 4332
rect 19628 3508 19648 4332
rect 18476 3480 19648 3508
rect 19888 4332 21060 4360
rect 19888 3508 20976 4332
rect 21040 3508 21060 4332
rect 19888 3480 21060 3508
rect 21300 4332 22472 4360
rect 21300 3508 22388 4332
rect 22452 3508 22472 4332
rect 21300 3480 22472 3508
rect 22712 4332 23884 4360
rect 22712 3508 23800 4332
rect 23864 3508 23884 4332
rect 22712 3480 23884 3508
rect -23884 3212 -22712 3240
rect -23884 2388 -22796 3212
rect -22732 2388 -22712 3212
rect -23884 2360 -22712 2388
rect -22472 3212 -21300 3240
rect -22472 2388 -21384 3212
rect -21320 2388 -21300 3212
rect -22472 2360 -21300 2388
rect -21060 3212 -19888 3240
rect -21060 2388 -19972 3212
rect -19908 2388 -19888 3212
rect -21060 2360 -19888 2388
rect -19648 3212 -18476 3240
rect -19648 2388 -18560 3212
rect -18496 2388 -18476 3212
rect -19648 2360 -18476 2388
rect -18236 3212 -17064 3240
rect -18236 2388 -17148 3212
rect -17084 2388 -17064 3212
rect -18236 2360 -17064 2388
rect -16824 3212 -15652 3240
rect -16824 2388 -15736 3212
rect -15672 2388 -15652 3212
rect -16824 2360 -15652 2388
rect -15412 3212 -14240 3240
rect -15412 2388 -14324 3212
rect -14260 2388 -14240 3212
rect -15412 2360 -14240 2388
rect -14000 3212 -12828 3240
rect -14000 2388 -12912 3212
rect -12848 2388 -12828 3212
rect -14000 2360 -12828 2388
rect -12588 3212 -11416 3240
rect -12588 2388 -11500 3212
rect -11436 2388 -11416 3212
rect -12588 2360 -11416 2388
rect -11176 3212 -10004 3240
rect -11176 2388 -10088 3212
rect -10024 2388 -10004 3212
rect -11176 2360 -10004 2388
rect -9764 3212 -8592 3240
rect -9764 2388 -8676 3212
rect -8612 2388 -8592 3212
rect -9764 2360 -8592 2388
rect -8352 3212 -7180 3240
rect -8352 2388 -7264 3212
rect -7200 2388 -7180 3212
rect -8352 2360 -7180 2388
rect -6940 3212 -5768 3240
rect -6940 2388 -5852 3212
rect -5788 2388 -5768 3212
rect -6940 2360 -5768 2388
rect -5528 3212 -4356 3240
rect -5528 2388 -4440 3212
rect -4376 2388 -4356 3212
rect -5528 2360 -4356 2388
rect -4116 3212 -2944 3240
rect -4116 2388 -3028 3212
rect -2964 2388 -2944 3212
rect -4116 2360 -2944 2388
rect -2704 3212 -1532 3240
rect -2704 2388 -1616 3212
rect -1552 2388 -1532 3212
rect -2704 2360 -1532 2388
rect -1292 3212 -120 3240
rect -1292 2388 -204 3212
rect -140 2388 -120 3212
rect -1292 2360 -120 2388
rect 120 3212 1292 3240
rect 120 2388 1208 3212
rect 1272 2388 1292 3212
rect 120 2360 1292 2388
rect 1532 3212 2704 3240
rect 1532 2388 2620 3212
rect 2684 2388 2704 3212
rect 1532 2360 2704 2388
rect 2944 3212 4116 3240
rect 2944 2388 4032 3212
rect 4096 2388 4116 3212
rect 2944 2360 4116 2388
rect 4356 3212 5528 3240
rect 4356 2388 5444 3212
rect 5508 2388 5528 3212
rect 4356 2360 5528 2388
rect 5768 3212 6940 3240
rect 5768 2388 6856 3212
rect 6920 2388 6940 3212
rect 5768 2360 6940 2388
rect 7180 3212 8352 3240
rect 7180 2388 8268 3212
rect 8332 2388 8352 3212
rect 7180 2360 8352 2388
rect 8592 3212 9764 3240
rect 8592 2388 9680 3212
rect 9744 2388 9764 3212
rect 8592 2360 9764 2388
rect 10004 3212 11176 3240
rect 10004 2388 11092 3212
rect 11156 2388 11176 3212
rect 10004 2360 11176 2388
rect 11416 3212 12588 3240
rect 11416 2388 12504 3212
rect 12568 2388 12588 3212
rect 11416 2360 12588 2388
rect 12828 3212 14000 3240
rect 12828 2388 13916 3212
rect 13980 2388 14000 3212
rect 12828 2360 14000 2388
rect 14240 3212 15412 3240
rect 14240 2388 15328 3212
rect 15392 2388 15412 3212
rect 14240 2360 15412 2388
rect 15652 3212 16824 3240
rect 15652 2388 16740 3212
rect 16804 2388 16824 3212
rect 15652 2360 16824 2388
rect 17064 3212 18236 3240
rect 17064 2388 18152 3212
rect 18216 2388 18236 3212
rect 17064 2360 18236 2388
rect 18476 3212 19648 3240
rect 18476 2388 19564 3212
rect 19628 2388 19648 3212
rect 18476 2360 19648 2388
rect 19888 3212 21060 3240
rect 19888 2388 20976 3212
rect 21040 2388 21060 3212
rect 19888 2360 21060 2388
rect 21300 3212 22472 3240
rect 21300 2388 22388 3212
rect 22452 2388 22472 3212
rect 21300 2360 22472 2388
rect 22712 3212 23884 3240
rect 22712 2388 23800 3212
rect 23864 2388 23884 3212
rect 22712 2360 23884 2388
rect -23884 2092 -22712 2120
rect -23884 1268 -22796 2092
rect -22732 1268 -22712 2092
rect -23884 1240 -22712 1268
rect -22472 2092 -21300 2120
rect -22472 1268 -21384 2092
rect -21320 1268 -21300 2092
rect -22472 1240 -21300 1268
rect -21060 2092 -19888 2120
rect -21060 1268 -19972 2092
rect -19908 1268 -19888 2092
rect -21060 1240 -19888 1268
rect -19648 2092 -18476 2120
rect -19648 1268 -18560 2092
rect -18496 1268 -18476 2092
rect -19648 1240 -18476 1268
rect -18236 2092 -17064 2120
rect -18236 1268 -17148 2092
rect -17084 1268 -17064 2092
rect -18236 1240 -17064 1268
rect -16824 2092 -15652 2120
rect -16824 1268 -15736 2092
rect -15672 1268 -15652 2092
rect -16824 1240 -15652 1268
rect -15412 2092 -14240 2120
rect -15412 1268 -14324 2092
rect -14260 1268 -14240 2092
rect -15412 1240 -14240 1268
rect -14000 2092 -12828 2120
rect -14000 1268 -12912 2092
rect -12848 1268 -12828 2092
rect -14000 1240 -12828 1268
rect -12588 2092 -11416 2120
rect -12588 1268 -11500 2092
rect -11436 1268 -11416 2092
rect -12588 1240 -11416 1268
rect -11176 2092 -10004 2120
rect -11176 1268 -10088 2092
rect -10024 1268 -10004 2092
rect -11176 1240 -10004 1268
rect -9764 2092 -8592 2120
rect -9764 1268 -8676 2092
rect -8612 1268 -8592 2092
rect -9764 1240 -8592 1268
rect -8352 2092 -7180 2120
rect -8352 1268 -7264 2092
rect -7200 1268 -7180 2092
rect -8352 1240 -7180 1268
rect -6940 2092 -5768 2120
rect -6940 1268 -5852 2092
rect -5788 1268 -5768 2092
rect -6940 1240 -5768 1268
rect -5528 2092 -4356 2120
rect -5528 1268 -4440 2092
rect -4376 1268 -4356 2092
rect -5528 1240 -4356 1268
rect -4116 2092 -2944 2120
rect -4116 1268 -3028 2092
rect -2964 1268 -2944 2092
rect -4116 1240 -2944 1268
rect -2704 2092 -1532 2120
rect -2704 1268 -1616 2092
rect -1552 1268 -1532 2092
rect -2704 1240 -1532 1268
rect -1292 2092 -120 2120
rect -1292 1268 -204 2092
rect -140 1268 -120 2092
rect -1292 1240 -120 1268
rect 120 2092 1292 2120
rect 120 1268 1208 2092
rect 1272 1268 1292 2092
rect 120 1240 1292 1268
rect 1532 2092 2704 2120
rect 1532 1268 2620 2092
rect 2684 1268 2704 2092
rect 1532 1240 2704 1268
rect 2944 2092 4116 2120
rect 2944 1268 4032 2092
rect 4096 1268 4116 2092
rect 2944 1240 4116 1268
rect 4356 2092 5528 2120
rect 4356 1268 5444 2092
rect 5508 1268 5528 2092
rect 4356 1240 5528 1268
rect 5768 2092 6940 2120
rect 5768 1268 6856 2092
rect 6920 1268 6940 2092
rect 5768 1240 6940 1268
rect 7180 2092 8352 2120
rect 7180 1268 8268 2092
rect 8332 1268 8352 2092
rect 7180 1240 8352 1268
rect 8592 2092 9764 2120
rect 8592 1268 9680 2092
rect 9744 1268 9764 2092
rect 8592 1240 9764 1268
rect 10004 2092 11176 2120
rect 10004 1268 11092 2092
rect 11156 1268 11176 2092
rect 10004 1240 11176 1268
rect 11416 2092 12588 2120
rect 11416 1268 12504 2092
rect 12568 1268 12588 2092
rect 11416 1240 12588 1268
rect 12828 2092 14000 2120
rect 12828 1268 13916 2092
rect 13980 1268 14000 2092
rect 12828 1240 14000 1268
rect 14240 2092 15412 2120
rect 14240 1268 15328 2092
rect 15392 1268 15412 2092
rect 14240 1240 15412 1268
rect 15652 2092 16824 2120
rect 15652 1268 16740 2092
rect 16804 1268 16824 2092
rect 15652 1240 16824 1268
rect 17064 2092 18236 2120
rect 17064 1268 18152 2092
rect 18216 1268 18236 2092
rect 17064 1240 18236 1268
rect 18476 2092 19648 2120
rect 18476 1268 19564 2092
rect 19628 1268 19648 2092
rect 18476 1240 19648 1268
rect 19888 2092 21060 2120
rect 19888 1268 20976 2092
rect 21040 1268 21060 2092
rect 19888 1240 21060 1268
rect 21300 2092 22472 2120
rect 21300 1268 22388 2092
rect 22452 1268 22472 2092
rect 21300 1240 22472 1268
rect 22712 2092 23884 2120
rect 22712 1268 23800 2092
rect 23864 1268 23884 2092
rect 22712 1240 23884 1268
rect -23884 972 -22712 1000
rect -23884 148 -22796 972
rect -22732 148 -22712 972
rect -23884 120 -22712 148
rect -22472 972 -21300 1000
rect -22472 148 -21384 972
rect -21320 148 -21300 972
rect -22472 120 -21300 148
rect -21060 972 -19888 1000
rect -21060 148 -19972 972
rect -19908 148 -19888 972
rect -21060 120 -19888 148
rect -19648 972 -18476 1000
rect -19648 148 -18560 972
rect -18496 148 -18476 972
rect -19648 120 -18476 148
rect -18236 972 -17064 1000
rect -18236 148 -17148 972
rect -17084 148 -17064 972
rect -18236 120 -17064 148
rect -16824 972 -15652 1000
rect -16824 148 -15736 972
rect -15672 148 -15652 972
rect -16824 120 -15652 148
rect -15412 972 -14240 1000
rect -15412 148 -14324 972
rect -14260 148 -14240 972
rect -15412 120 -14240 148
rect -14000 972 -12828 1000
rect -14000 148 -12912 972
rect -12848 148 -12828 972
rect -14000 120 -12828 148
rect -12588 972 -11416 1000
rect -12588 148 -11500 972
rect -11436 148 -11416 972
rect -12588 120 -11416 148
rect -11176 972 -10004 1000
rect -11176 148 -10088 972
rect -10024 148 -10004 972
rect -11176 120 -10004 148
rect -9764 972 -8592 1000
rect -9764 148 -8676 972
rect -8612 148 -8592 972
rect -9764 120 -8592 148
rect -8352 972 -7180 1000
rect -8352 148 -7264 972
rect -7200 148 -7180 972
rect -8352 120 -7180 148
rect -6940 972 -5768 1000
rect -6940 148 -5852 972
rect -5788 148 -5768 972
rect -6940 120 -5768 148
rect -5528 972 -4356 1000
rect -5528 148 -4440 972
rect -4376 148 -4356 972
rect -5528 120 -4356 148
rect -4116 972 -2944 1000
rect -4116 148 -3028 972
rect -2964 148 -2944 972
rect -4116 120 -2944 148
rect -2704 972 -1532 1000
rect -2704 148 -1616 972
rect -1552 148 -1532 972
rect -2704 120 -1532 148
rect -1292 972 -120 1000
rect -1292 148 -204 972
rect -140 148 -120 972
rect -1292 120 -120 148
rect 120 972 1292 1000
rect 120 148 1208 972
rect 1272 148 1292 972
rect 120 120 1292 148
rect 1532 972 2704 1000
rect 1532 148 2620 972
rect 2684 148 2704 972
rect 1532 120 2704 148
rect 2944 972 4116 1000
rect 2944 148 4032 972
rect 4096 148 4116 972
rect 2944 120 4116 148
rect 4356 972 5528 1000
rect 4356 148 5444 972
rect 5508 148 5528 972
rect 4356 120 5528 148
rect 5768 972 6940 1000
rect 5768 148 6856 972
rect 6920 148 6940 972
rect 5768 120 6940 148
rect 7180 972 8352 1000
rect 7180 148 8268 972
rect 8332 148 8352 972
rect 7180 120 8352 148
rect 8592 972 9764 1000
rect 8592 148 9680 972
rect 9744 148 9764 972
rect 8592 120 9764 148
rect 10004 972 11176 1000
rect 10004 148 11092 972
rect 11156 148 11176 972
rect 10004 120 11176 148
rect 11416 972 12588 1000
rect 11416 148 12504 972
rect 12568 148 12588 972
rect 11416 120 12588 148
rect 12828 972 14000 1000
rect 12828 148 13916 972
rect 13980 148 14000 972
rect 12828 120 14000 148
rect 14240 972 15412 1000
rect 14240 148 15328 972
rect 15392 148 15412 972
rect 14240 120 15412 148
rect 15652 972 16824 1000
rect 15652 148 16740 972
rect 16804 148 16824 972
rect 15652 120 16824 148
rect 17064 972 18236 1000
rect 17064 148 18152 972
rect 18216 148 18236 972
rect 17064 120 18236 148
rect 18476 972 19648 1000
rect 18476 148 19564 972
rect 19628 148 19648 972
rect 18476 120 19648 148
rect 19888 972 21060 1000
rect 19888 148 20976 972
rect 21040 148 21060 972
rect 19888 120 21060 148
rect 21300 972 22472 1000
rect 21300 148 22388 972
rect 22452 148 22472 972
rect 21300 120 22472 148
rect 22712 972 23884 1000
rect 22712 148 23800 972
rect 23864 148 23884 972
rect 22712 120 23884 148
rect -23884 -148 -22712 -120
rect -23884 -972 -22796 -148
rect -22732 -972 -22712 -148
rect -23884 -1000 -22712 -972
rect -22472 -148 -21300 -120
rect -22472 -972 -21384 -148
rect -21320 -972 -21300 -148
rect -22472 -1000 -21300 -972
rect -21060 -148 -19888 -120
rect -21060 -972 -19972 -148
rect -19908 -972 -19888 -148
rect -21060 -1000 -19888 -972
rect -19648 -148 -18476 -120
rect -19648 -972 -18560 -148
rect -18496 -972 -18476 -148
rect -19648 -1000 -18476 -972
rect -18236 -148 -17064 -120
rect -18236 -972 -17148 -148
rect -17084 -972 -17064 -148
rect -18236 -1000 -17064 -972
rect -16824 -148 -15652 -120
rect -16824 -972 -15736 -148
rect -15672 -972 -15652 -148
rect -16824 -1000 -15652 -972
rect -15412 -148 -14240 -120
rect -15412 -972 -14324 -148
rect -14260 -972 -14240 -148
rect -15412 -1000 -14240 -972
rect -14000 -148 -12828 -120
rect -14000 -972 -12912 -148
rect -12848 -972 -12828 -148
rect -14000 -1000 -12828 -972
rect -12588 -148 -11416 -120
rect -12588 -972 -11500 -148
rect -11436 -972 -11416 -148
rect -12588 -1000 -11416 -972
rect -11176 -148 -10004 -120
rect -11176 -972 -10088 -148
rect -10024 -972 -10004 -148
rect -11176 -1000 -10004 -972
rect -9764 -148 -8592 -120
rect -9764 -972 -8676 -148
rect -8612 -972 -8592 -148
rect -9764 -1000 -8592 -972
rect -8352 -148 -7180 -120
rect -8352 -972 -7264 -148
rect -7200 -972 -7180 -148
rect -8352 -1000 -7180 -972
rect -6940 -148 -5768 -120
rect -6940 -972 -5852 -148
rect -5788 -972 -5768 -148
rect -6940 -1000 -5768 -972
rect -5528 -148 -4356 -120
rect -5528 -972 -4440 -148
rect -4376 -972 -4356 -148
rect -5528 -1000 -4356 -972
rect -4116 -148 -2944 -120
rect -4116 -972 -3028 -148
rect -2964 -972 -2944 -148
rect -4116 -1000 -2944 -972
rect -2704 -148 -1532 -120
rect -2704 -972 -1616 -148
rect -1552 -972 -1532 -148
rect -2704 -1000 -1532 -972
rect -1292 -148 -120 -120
rect -1292 -972 -204 -148
rect -140 -972 -120 -148
rect -1292 -1000 -120 -972
rect 120 -148 1292 -120
rect 120 -972 1208 -148
rect 1272 -972 1292 -148
rect 120 -1000 1292 -972
rect 1532 -148 2704 -120
rect 1532 -972 2620 -148
rect 2684 -972 2704 -148
rect 1532 -1000 2704 -972
rect 2944 -148 4116 -120
rect 2944 -972 4032 -148
rect 4096 -972 4116 -148
rect 2944 -1000 4116 -972
rect 4356 -148 5528 -120
rect 4356 -972 5444 -148
rect 5508 -972 5528 -148
rect 4356 -1000 5528 -972
rect 5768 -148 6940 -120
rect 5768 -972 6856 -148
rect 6920 -972 6940 -148
rect 5768 -1000 6940 -972
rect 7180 -148 8352 -120
rect 7180 -972 8268 -148
rect 8332 -972 8352 -148
rect 7180 -1000 8352 -972
rect 8592 -148 9764 -120
rect 8592 -972 9680 -148
rect 9744 -972 9764 -148
rect 8592 -1000 9764 -972
rect 10004 -148 11176 -120
rect 10004 -972 11092 -148
rect 11156 -972 11176 -148
rect 10004 -1000 11176 -972
rect 11416 -148 12588 -120
rect 11416 -972 12504 -148
rect 12568 -972 12588 -148
rect 11416 -1000 12588 -972
rect 12828 -148 14000 -120
rect 12828 -972 13916 -148
rect 13980 -972 14000 -148
rect 12828 -1000 14000 -972
rect 14240 -148 15412 -120
rect 14240 -972 15328 -148
rect 15392 -972 15412 -148
rect 14240 -1000 15412 -972
rect 15652 -148 16824 -120
rect 15652 -972 16740 -148
rect 16804 -972 16824 -148
rect 15652 -1000 16824 -972
rect 17064 -148 18236 -120
rect 17064 -972 18152 -148
rect 18216 -972 18236 -148
rect 17064 -1000 18236 -972
rect 18476 -148 19648 -120
rect 18476 -972 19564 -148
rect 19628 -972 19648 -148
rect 18476 -1000 19648 -972
rect 19888 -148 21060 -120
rect 19888 -972 20976 -148
rect 21040 -972 21060 -148
rect 19888 -1000 21060 -972
rect 21300 -148 22472 -120
rect 21300 -972 22388 -148
rect 22452 -972 22472 -148
rect 21300 -1000 22472 -972
rect 22712 -148 23884 -120
rect 22712 -972 23800 -148
rect 23864 -972 23884 -148
rect 22712 -1000 23884 -972
rect -23884 -1268 -22712 -1240
rect -23884 -2092 -22796 -1268
rect -22732 -2092 -22712 -1268
rect -23884 -2120 -22712 -2092
rect -22472 -1268 -21300 -1240
rect -22472 -2092 -21384 -1268
rect -21320 -2092 -21300 -1268
rect -22472 -2120 -21300 -2092
rect -21060 -1268 -19888 -1240
rect -21060 -2092 -19972 -1268
rect -19908 -2092 -19888 -1268
rect -21060 -2120 -19888 -2092
rect -19648 -1268 -18476 -1240
rect -19648 -2092 -18560 -1268
rect -18496 -2092 -18476 -1268
rect -19648 -2120 -18476 -2092
rect -18236 -1268 -17064 -1240
rect -18236 -2092 -17148 -1268
rect -17084 -2092 -17064 -1268
rect -18236 -2120 -17064 -2092
rect -16824 -1268 -15652 -1240
rect -16824 -2092 -15736 -1268
rect -15672 -2092 -15652 -1268
rect -16824 -2120 -15652 -2092
rect -15412 -1268 -14240 -1240
rect -15412 -2092 -14324 -1268
rect -14260 -2092 -14240 -1268
rect -15412 -2120 -14240 -2092
rect -14000 -1268 -12828 -1240
rect -14000 -2092 -12912 -1268
rect -12848 -2092 -12828 -1268
rect -14000 -2120 -12828 -2092
rect -12588 -1268 -11416 -1240
rect -12588 -2092 -11500 -1268
rect -11436 -2092 -11416 -1268
rect -12588 -2120 -11416 -2092
rect -11176 -1268 -10004 -1240
rect -11176 -2092 -10088 -1268
rect -10024 -2092 -10004 -1268
rect -11176 -2120 -10004 -2092
rect -9764 -1268 -8592 -1240
rect -9764 -2092 -8676 -1268
rect -8612 -2092 -8592 -1268
rect -9764 -2120 -8592 -2092
rect -8352 -1268 -7180 -1240
rect -8352 -2092 -7264 -1268
rect -7200 -2092 -7180 -1268
rect -8352 -2120 -7180 -2092
rect -6940 -1268 -5768 -1240
rect -6940 -2092 -5852 -1268
rect -5788 -2092 -5768 -1268
rect -6940 -2120 -5768 -2092
rect -5528 -1268 -4356 -1240
rect -5528 -2092 -4440 -1268
rect -4376 -2092 -4356 -1268
rect -5528 -2120 -4356 -2092
rect -4116 -1268 -2944 -1240
rect -4116 -2092 -3028 -1268
rect -2964 -2092 -2944 -1268
rect -4116 -2120 -2944 -2092
rect -2704 -1268 -1532 -1240
rect -2704 -2092 -1616 -1268
rect -1552 -2092 -1532 -1268
rect -2704 -2120 -1532 -2092
rect -1292 -1268 -120 -1240
rect -1292 -2092 -204 -1268
rect -140 -2092 -120 -1268
rect -1292 -2120 -120 -2092
rect 120 -1268 1292 -1240
rect 120 -2092 1208 -1268
rect 1272 -2092 1292 -1268
rect 120 -2120 1292 -2092
rect 1532 -1268 2704 -1240
rect 1532 -2092 2620 -1268
rect 2684 -2092 2704 -1268
rect 1532 -2120 2704 -2092
rect 2944 -1268 4116 -1240
rect 2944 -2092 4032 -1268
rect 4096 -2092 4116 -1268
rect 2944 -2120 4116 -2092
rect 4356 -1268 5528 -1240
rect 4356 -2092 5444 -1268
rect 5508 -2092 5528 -1268
rect 4356 -2120 5528 -2092
rect 5768 -1268 6940 -1240
rect 5768 -2092 6856 -1268
rect 6920 -2092 6940 -1268
rect 5768 -2120 6940 -2092
rect 7180 -1268 8352 -1240
rect 7180 -2092 8268 -1268
rect 8332 -2092 8352 -1268
rect 7180 -2120 8352 -2092
rect 8592 -1268 9764 -1240
rect 8592 -2092 9680 -1268
rect 9744 -2092 9764 -1268
rect 8592 -2120 9764 -2092
rect 10004 -1268 11176 -1240
rect 10004 -2092 11092 -1268
rect 11156 -2092 11176 -1268
rect 10004 -2120 11176 -2092
rect 11416 -1268 12588 -1240
rect 11416 -2092 12504 -1268
rect 12568 -2092 12588 -1268
rect 11416 -2120 12588 -2092
rect 12828 -1268 14000 -1240
rect 12828 -2092 13916 -1268
rect 13980 -2092 14000 -1268
rect 12828 -2120 14000 -2092
rect 14240 -1268 15412 -1240
rect 14240 -2092 15328 -1268
rect 15392 -2092 15412 -1268
rect 14240 -2120 15412 -2092
rect 15652 -1268 16824 -1240
rect 15652 -2092 16740 -1268
rect 16804 -2092 16824 -1268
rect 15652 -2120 16824 -2092
rect 17064 -1268 18236 -1240
rect 17064 -2092 18152 -1268
rect 18216 -2092 18236 -1268
rect 17064 -2120 18236 -2092
rect 18476 -1268 19648 -1240
rect 18476 -2092 19564 -1268
rect 19628 -2092 19648 -1268
rect 18476 -2120 19648 -2092
rect 19888 -1268 21060 -1240
rect 19888 -2092 20976 -1268
rect 21040 -2092 21060 -1268
rect 19888 -2120 21060 -2092
rect 21300 -1268 22472 -1240
rect 21300 -2092 22388 -1268
rect 22452 -2092 22472 -1268
rect 21300 -2120 22472 -2092
rect 22712 -1268 23884 -1240
rect 22712 -2092 23800 -1268
rect 23864 -2092 23884 -1268
rect 22712 -2120 23884 -2092
rect -23884 -2388 -22712 -2360
rect -23884 -3212 -22796 -2388
rect -22732 -3212 -22712 -2388
rect -23884 -3240 -22712 -3212
rect -22472 -2388 -21300 -2360
rect -22472 -3212 -21384 -2388
rect -21320 -3212 -21300 -2388
rect -22472 -3240 -21300 -3212
rect -21060 -2388 -19888 -2360
rect -21060 -3212 -19972 -2388
rect -19908 -3212 -19888 -2388
rect -21060 -3240 -19888 -3212
rect -19648 -2388 -18476 -2360
rect -19648 -3212 -18560 -2388
rect -18496 -3212 -18476 -2388
rect -19648 -3240 -18476 -3212
rect -18236 -2388 -17064 -2360
rect -18236 -3212 -17148 -2388
rect -17084 -3212 -17064 -2388
rect -18236 -3240 -17064 -3212
rect -16824 -2388 -15652 -2360
rect -16824 -3212 -15736 -2388
rect -15672 -3212 -15652 -2388
rect -16824 -3240 -15652 -3212
rect -15412 -2388 -14240 -2360
rect -15412 -3212 -14324 -2388
rect -14260 -3212 -14240 -2388
rect -15412 -3240 -14240 -3212
rect -14000 -2388 -12828 -2360
rect -14000 -3212 -12912 -2388
rect -12848 -3212 -12828 -2388
rect -14000 -3240 -12828 -3212
rect -12588 -2388 -11416 -2360
rect -12588 -3212 -11500 -2388
rect -11436 -3212 -11416 -2388
rect -12588 -3240 -11416 -3212
rect -11176 -2388 -10004 -2360
rect -11176 -3212 -10088 -2388
rect -10024 -3212 -10004 -2388
rect -11176 -3240 -10004 -3212
rect -9764 -2388 -8592 -2360
rect -9764 -3212 -8676 -2388
rect -8612 -3212 -8592 -2388
rect -9764 -3240 -8592 -3212
rect -8352 -2388 -7180 -2360
rect -8352 -3212 -7264 -2388
rect -7200 -3212 -7180 -2388
rect -8352 -3240 -7180 -3212
rect -6940 -2388 -5768 -2360
rect -6940 -3212 -5852 -2388
rect -5788 -3212 -5768 -2388
rect -6940 -3240 -5768 -3212
rect -5528 -2388 -4356 -2360
rect -5528 -3212 -4440 -2388
rect -4376 -3212 -4356 -2388
rect -5528 -3240 -4356 -3212
rect -4116 -2388 -2944 -2360
rect -4116 -3212 -3028 -2388
rect -2964 -3212 -2944 -2388
rect -4116 -3240 -2944 -3212
rect -2704 -2388 -1532 -2360
rect -2704 -3212 -1616 -2388
rect -1552 -3212 -1532 -2388
rect -2704 -3240 -1532 -3212
rect -1292 -2388 -120 -2360
rect -1292 -3212 -204 -2388
rect -140 -3212 -120 -2388
rect -1292 -3240 -120 -3212
rect 120 -2388 1292 -2360
rect 120 -3212 1208 -2388
rect 1272 -3212 1292 -2388
rect 120 -3240 1292 -3212
rect 1532 -2388 2704 -2360
rect 1532 -3212 2620 -2388
rect 2684 -3212 2704 -2388
rect 1532 -3240 2704 -3212
rect 2944 -2388 4116 -2360
rect 2944 -3212 4032 -2388
rect 4096 -3212 4116 -2388
rect 2944 -3240 4116 -3212
rect 4356 -2388 5528 -2360
rect 4356 -3212 5444 -2388
rect 5508 -3212 5528 -2388
rect 4356 -3240 5528 -3212
rect 5768 -2388 6940 -2360
rect 5768 -3212 6856 -2388
rect 6920 -3212 6940 -2388
rect 5768 -3240 6940 -3212
rect 7180 -2388 8352 -2360
rect 7180 -3212 8268 -2388
rect 8332 -3212 8352 -2388
rect 7180 -3240 8352 -3212
rect 8592 -2388 9764 -2360
rect 8592 -3212 9680 -2388
rect 9744 -3212 9764 -2388
rect 8592 -3240 9764 -3212
rect 10004 -2388 11176 -2360
rect 10004 -3212 11092 -2388
rect 11156 -3212 11176 -2388
rect 10004 -3240 11176 -3212
rect 11416 -2388 12588 -2360
rect 11416 -3212 12504 -2388
rect 12568 -3212 12588 -2388
rect 11416 -3240 12588 -3212
rect 12828 -2388 14000 -2360
rect 12828 -3212 13916 -2388
rect 13980 -3212 14000 -2388
rect 12828 -3240 14000 -3212
rect 14240 -2388 15412 -2360
rect 14240 -3212 15328 -2388
rect 15392 -3212 15412 -2388
rect 14240 -3240 15412 -3212
rect 15652 -2388 16824 -2360
rect 15652 -3212 16740 -2388
rect 16804 -3212 16824 -2388
rect 15652 -3240 16824 -3212
rect 17064 -2388 18236 -2360
rect 17064 -3212 18152 -2388
rect 18216 -3212 18236 -2388
rect 17064 -3240 18236 -3212
rect 18476 -2388 19648 -2360
rect 18476 -3212 19564 -2388
rect 19628 -3212 19648 -2388
rect 18476 -3240 19648 -3212
rect 19888 -2388 21060 -2360
rect 19888 -3212 20976 -2388
rect 21040 -3212 21060 -2388
rect 19888 -3240 21060 -3212
rect 21300 -2388 22472 -2360
rect 21300 -3212 22388 -2388
rect 22452 -3212 22472 -2388
rect 21300 -3240 22472 -3212
rect 22712 -2388 23884 -2360
rect 22712 -3212 23800 -2388
rect 23864 -3212 23884 -2388
rect 22712 -3240 23884 -3212
rect -23884 -3508 -22712 -3480
rect -23884 -4332 -22796 -3508
rect -22732 -4332 -22712 -3508
rect -23884 -4360 -22712 -4332
rect -22472 -3508 -21300 -3480
rect -22472 -4332 -21384 -3508
rect -21320 -4332 -21300 -3508
rect -22472 -4360 -21300 -4332
rect -21060 -3508 -19888 -3480
rect -21060 -4332 -19972 -3508
rect -19908 -4332 -19888 -3508
rect -21060 -4360 -19888 -4332
rect -19648 -3508 -18476 -3480
rect -19648 -4332 -18560 -3508
rect -18496 -4332 -18476 -3508
rect -19648 -4360 -18476 -4332
rect -18236 -3508 -17064 -3480
rect -18236 -4332 -17148 -3508
rect -17084 -4332 -17064 -3508
rect -18236 -4360 -17064 -4332
rect -16824 -3508 -15652 -3480
rect -16824 -4332 -15736 -3508
rect -15672 -4332 -15652 -3508
rect -16824 -4360 -15652 -4332
rect -15412 -3508 -14240 -3480
rect -15412 -4332 -14324 -3508
rect -14260 -4332 -14240 -3508
rect -15412 -4360 -14240 -4332
rect -14000 -3508 -12828 -3480
rect -14000 -4332 -12912 -3508
rect -12848 -4332 -12828 -3508
rect -14000 -4360 -12828 -4332
rect -12588 -3508 -11416 -3480
rect -12588 -4332 -11500 -3508
rect -11436 -4332 -11416 -3508
rect -12588 -4360 -11416 -4332
rect -11176 -3508 -10004 -3480
rect -11176 -4332 -10088 -3508
rect -10024 -4332 -10004 -3508
rect -11176 -4360 -10004 -4332
rect -9764 -3508 -8592 -3480
rect -9764 -4332 -8676 -3508
rect -8612 -4332 -8592 -3508
rect -9764 -4360 -8592 -4332
rect -8352 -3508 -7180 -3480
rect -8352 -4332 -7264 -3508
rect -7200 -4332 -7180 -3508
rect -8352 -4360 -7180 -4332
rect -6940 -3508 -5768 -3480
rect -6940 -4332 -5852 -3508
rect -5788 -4332 -5768 -3508
rect -6940 -4360 -5768 -4332
rect -5528 -3508 -4356 -3480
rect -5528 -4332 -4440 -3508
rect -4376 -4332 -4356 -3508
rect -5528 -4360 -4356 -4332
rect -4116 -3508 -2944 -3480
rect -4116 -4332 -3028 -3508
rect -2964 -4332 -2944 -3508
rect -4116 -4360 -2944 -4332
rect -2704 -3508 -1532 -3480
rect -2704 -4332 -1616 -3508
rect -1552 -4332 -1532 -3508
rect -2704 -4360 -1532 -4332
rect -1292 -3508 -120 -3480
rect -1292 -4332 -204 -3508
rect -140 -4332 -120 -3508
rect -1292 -4360 -120 -4332
rect 120 -3508 1292 -3480
rect 120 -4332 1208 -3508
rect 1272 -4332 1292 -3508
rect 120 -4360 1292 -4332
rect 1532 -3508 2704 -3480
rect 1532 -4332 2620 -3508
rect 2684 -4332 2704 -3508
rect 1532 -4360 2704 -4332
rect 2944 -3508 4116 -3480
rect 2944 -4332 4032 -3508
rect 4096 -4332 4116 -3508
rect 2944 -4360 4116 -4332
rect 4356 -3508 5528 -3480
rect 4356 -4332 5444 -3508
rect 5508 -4332 5528 -3508
rect 4356 -4360 5528 -4332
rect 5768 -3508 6940 -3480
rect 5768 -4332 6856 -3508
rect 6920 -4332 6940 -3508
rect 5768 -4360 6940 -4332
rect 7180 -3508 8352 -3480
rect 7180 -4332 8268 -3508
rect 8332 -4332 8352 -3508
rect 7180 -4360 8352 -4332
rect 8592 -3508 9764 -3480
rect 8592 -4332 9680 -3508
rect 9744 -4332 9764 -3508
rect 8592 -4360 9764 -4332
rect 10004 -3508 11176 -3480
rect 10004 -4332 11092 -3508
rect 11156 -4332 11176 -3508
rect 10004 -4360 11176 -4332
rect 11416 -3508 12588 -3480
rect 11416 -4332 12504 -3508
rect 12568 -4332 12588 -3508
rect 11416 -4360 12588 -4332
rect 12828 -3508 14000 -3480
rect 12828 -4332 13916 -3508
rect 13980 -4332 14000 -3508
rect 12828 -4360 14000 -4332
rect 14240 -3508 15412 -3480
rect 14240 -4332 15328 -3508
rect 15392 -4332 15412 -3508
rect 14240 -4360 15412 -4332
rect 15652 -3508 16824 -3480
rect 15652 -4332 16740 -3508
rect 16804 -4332 16824 -3508
rect 15652 -4360 16824 -4332
rect 17064 -3508 18236 -3480
rect 17064 -4332 18152 -3508
rect 18216 -4332 18236 -3508
rect 17064 -4360 18236 -4332
rect 18476 -3508 19648 -3480
rect 18476 -4332 19564 -3508
rect 19628 -4332 19648 -3508
rect 18476 -4360 19648 -4332
rect 19888 -3508 21060 -3480
rect 19888 -4332 20976 -3508
rect 21040 -4332 21060 -3508
rect 19888 -4360 21060 -4332
rect 21300 -3508 22472 -3480
rect 21300 -4332 22388 -3508
rect 22452 -4332 22472 -3508
rect 21300 -4360 22472 -4332
rect 22712 -3508 23884 -3480
rect 22712 -4332 23800 -3508
rect 23864 -4332 23884 -3508
rect 22712 -4360 23884 -4332
rect -23884 -4628 -22712 -4600
rect -23884 -5452 -22796 -4628
rect -22732 -5452 -22712 -4628
rect -23884 -5480 -22712 -5452
rect -22472 -4628 -21300 -4600
rect -22472 -5452 -21384 -4628
rect -21320 -5452 -21300 -4628
rect -22472 -5480 -21300 -5452
rect -21060 -4628 -19888 -4600
rect -21060 -5452 -19972 -4628
rect -19908 -5452 -19888 -4628
rect -21060 -5480 -19888 -5452
rect -19648 -4628 -18476 -4600
rect -19648 -5452 -18560 -4628
rect -18496 -5452 -18476 -4628
rect -19648 -5480 -18476 -5452
rect -18236 -4628 -17064 -4600
rect -18236 -5452 -17148 -4628
rect -17084 -5452 -17064 -4628
rect -18236 -5480 -17064 -5452
rect -16824 -4628 -15652 -4600
rect -16824 -5452 -15736 -4628
rect -15672 -5452 -15652 -4628
rect -16824 -5480 -15652 -5452
rect -15412 -4628 -14240 -4600
rect -15412 -5452 -14324 -4628
rect -14260 -5452 -14240 -4628
rect -15412 -5480 -14240 -5452
rect -14000 -4628 -12828 -4600
rect -14000 -5452 -12912 -4628
rect -12848 -5452 -12828 -4628
rect -14000 -5480 -12828 -5452
rect -12588 -4628 -11416 -4600
rect -12588 -5452 -11500 -4628
rect -11436 -5452 -11416 -4628
rect -12588 -5480 -11416 -5452
rect -11176 -4628 -10004 -4600
rect -11176 -5452 -10088 -4628
rect -10024 -5452 -10004 -4628
rect -11176 -5480 -10004 -5452
rect -9764 -4628 -8592 -4600
rect -9764 -5452 -8676 -4628
rect -8612 -5452 -8592 -4628
rect -9764 -5480 -8592 -5452
rect -8352 -4628 -7180 -4600
rect -8352 -5452 -7264 -4628
rect -7200 -5452 -7180 -4628
rect -8352 -5480 -7180 -5452
rect -6940 -4628 -5768 -4600
rect -6940 -5452 -5852 -4628
rect -5788 -5452 -5768 -4628
rect -6940 -5480 -5768 -5452
rect -5528 -4628 -4356 -4600
rect -5528 -5452 -4440 -4628
rect -4376 -5452 -4356 -4628
rect -5528 -5480 -4356 -5452
rect -4116 -4628 -2944 -4600
rect -4116 -5452 -3028 -4628
rect -2964 -5452 -2944 -4628
rect -4116 -5480 -2944 -5452
rect -2704 -4628 -1532 -4600
rect -2704 -5452 -1616 -4628
rect -1552 -5452 -1532 -4628
rect -2704 -5480 -1532 -5452
rect -1292 -4628 -120 -4600
rect -1292 -5452 -204 -4628
rect -140 -5452 -120 -4628
rect -1292 -5480 -120 -5452
rect 120 -4628 1292 -4600
rect 120 -5452 1208 -4628
rect 1272 -5452 1292 -4628
rect 120 -5480 1292 -5452
rect 1532 -4628 2704 -4600
rect 1532 -5452 2620 -4628
rect 2684 -5452 2704 -4628
rect 1532 -5480 2704 -5452
rect 2944 -4628 4116 -4600
rect 2944 -5452 4032 -4628
rect 4096 -5452 4116 -4628
rect 2944 -5480 4116 -5452
rect 4356 -4628 5528 -4600
rect 4356 -5452 5444 -4628
rect 5508 -5452 5528 -4628
rect 4356 -5480 5528 -5452
rect 5768 -4628 6940 -4600
rect 5768 -5452 6856 -4628
rect 6920 -5452 6940 -4628
rect 5768 -5480 6940 -5452
rect 7180 -4628 8352 -4600
rect 7180 -5452 8268 -4628
rect 8332 -5452 8352 -4628
rect 7180 -5480 8352 -5452
rect 8592 -4628 9764 -4600
rect 8592 -5452 9680 -4628
rect 9744 -5452 9764 -4628
rect 8592 -5480 9764 -5452
rect 10004 -4628 11176 -4600
rect 10004 -5452 11092 -4628
rect 11156 -5452 11176 -4628
rect 10004 -5480 11176 -5452
rect 11416 -4628 12588 -4600
rect 11416 -5452 12504 -4628
rect 12568 -5452 12588 -4628
rect 11416 -5480 12588 -5452
rect 12828 -4628 14000 -4600
rect 12828 -5452 13916 -4628
rect 13980 -5452 14000 -4628
rect 12828 -5480 14000 -5452
rect 14240 -4628 15412 -4600
rect 14240 -5452 15328 -4628
rect 15392 -5452 15412 -4628
rect 14240 -5480 15412 -5452
rect 15652 -4628 16824 -4600
rect 15652 -5452 16740 -4628
rect 16804 -5452 16824 -4628
rect 15652 -5480 16824 -5452
rect 17064 -4628 18236 -4600
rect 17064 -5452 18152 -4628
rect 18216 -5452 18236 -4628
rect 17064 -5480 18236 -5452
rect 18476 -4628 19648 -4600
rect 18476 -5452 19564 -4628
rect 19628 -5452 19648 -4628
rect 18476 -5480 19648 -5452
rect 19888 -4628 21060 -4600
rect 19888 -5452 20976 -4628
rect 21040 -5452 21060 -4628
rect 19888 -5480 21060 -5452
rect 21300 -4628 22472 -4600
rect 21300 -5452 22388 -4628
rect 22452 -5452 22472 -4628
rect 21300 -5480 22472 -5452
rect 22712 -4628 23884 -4600
rect 22712 -5452 23800 -4628
rect 23864 -5452 23884 -4628
rect 22712 -5480 23884 -5452
rect -23884 -5748 -22712 -5720
rect -23884 -6572 -22796 -5748
rect -22732 -6572 -22712 -5748
rect -23884 -6600 -22712 -6572
rect -22472 -5748 -21300 -5720
rect -22472 -6572 -21384 -5748
rect -21320 -6572 -21300 -5748
rect -22472 -6600 -21300 -6572
rect -21060 -5748 -19888 -5720
rect -21060 -6572 -19972 -5748
rect -19908 -6572 -19888 -5748
rect -21060 -6600 -19888 -6572
rect -19648 -5748 -18476 -5720
rect -19648 -6572 -18560 -5748
rect -18496 -6572 -18476 -5748
rect -19648 -6600 -18476 -6572
rect -18236 -5748 -17064 -5720
rect -18236 -6572 -17148 -5748
rect -17084 -6572 -17064 -5748
rect -18236 -6600 -17064 -6572
rect -16824 -5748 -15652 -5720
rect -16824 -6572 -15736 -5748
rect -15672 -6572 -15652 -5748
rect -16824 -6600 -15652 -6572
rect -15412 -5748 -14240 -5720
rect -15412 -6572 -14324 -5748
rect -14260 -6572 -14240 -5748
rect -15412 -6600 -14240 -6572
rect -14000 -5748 -12828 -5720
rect -14000 -6572 -12912 -5748
rect -12848 -6572 -12828 -5748
rect -14000 -6600 -12828 -6572
rect -12588 -5748 -11416 -5720
rect -12588 -6572 -11500 -5748
rect -11436 -6572 -11416 -5748
rect -12588 -6600 -11416 -6572
rect -11176 -5748 -10004 -5720
rect -11176 -6572 -10088 -5748
rect -10024 -6572 -10004 -5748
rect -11176 -6600 -10004 -6572
rect -9764 -5748 -8592 -5720
rect -9764 -6572 -8676 -5748
rect -8612 -6572 -8592 -5748
rect -9764 -6600 -8592 -6572
rect -8352 -5748 -7180 -5720
rect -8352 -6572 -7264 -5748
rect -7200 -6572 -7180 -5748
rect -8352 -6600 -7180 -6572
rect -6940 -5748 -5768 -5720
rect -6940 -6572 -5852 -5748
rect -5788 -6572 -5768 -5748
rect -6940 -6600 -5768 -6572
rect -5528 -5748 -4356 -5720
rect -5528 -6572 -4440 -5748
rect -4376 -6572 -4356 -5748
rect -5528 -6600 -4356 -6572
rect -4116 -5748 -2944 -5720
rect -4116 -6572 -3028 -5748
rect -2964 -6572 -2944 -5748
rect -4116 -6600 -2944 -6572
rect -2704 -5748 -1532 -5720
rect -2704 -6572 -1616 -5748
rect -1552 -6572 -1532 -5748
rect -2704 -6600 -1532 -6572
rect -1292 -5748 -120 -5720
rect -1292 -6572 -204 -5748
rect -140 -6572 -120 -5748
rect -1292 -6600 -120 -6572
rect 120 -5748 1292 -5720
rect 120 -6572 1208 -5748
rect 1272 -6572 1292 -5748
rect 120 -6600 1292 -6572
rect 1532 -5748 2704 -5720
rect 1532 -6572 2620 -5748
rect 2684 -6572 2704 -5748
rect 1532 -6600 2704 -6572
rect 2944 -5748 4116 -5720
rect 2944 -6572 4032 -5748
rect 4096 -6572 4116 -5748
rect 2944 -6600 4116 -6572
rect 4356 -5748 5528 -5720
rect 4356 -6572 5444 -5748
rect 5508 -6572 5528 -5748
rect 4356 -6600 5528 -6572
rect 5768 -5748 6940 -5720
rect 5768 -6572 6856 -5748
rect 6920 -6572 6940 -5748
rect 5768 -6600 6940 -6572
rect 7180 -5748 8352 -5720
rect 7180 -6572 8268 -5748
rect 8332 -6572 8352 -5748
rect 7180 -6600 8352 -6572
rect 8592 -5748 9764 -5720
rect 8592 -6572 9680 -5748
rect 9744 -6572 9764 -5748
rect 8592 -6600 9764 -6572
rect 10004 -5748 11176 -5720
rect 10004 -6572 11092 -5748
rect 11156 -6572 11176 -5748
rect 10004 -6600 11176 -6572
rect 11416 -5748 12588 -5720
rect 11416 -6572 12504 -5748
rect 12568 -6572 12588 -5748
rect 11416 -6600 12588 -6572
rect 12828 -5748 14000 -5720
rect 12828 -6572 13916 -5748
rect 13980 -6572 14000 -5748
rect 12828 -6600 14000 -6572
rect 14240 -5748 15412 -5720
rect 14240 -6572 15328 -5748
rect 15392 -6572 15412 -5748
rect 14240 -6600 15412 -6572
rect 15652 -5748 16824 -5720
rect 15652 -6572 16740 -5748
rect 16804 -6572 16824 -5748
rect 15652 -6600 16824 -6572
rect 17064 -5748 18236 -5720
rect 17064 -6572 18152 -5748
rect 18216 -6572 18236 -5748
rect 17064 -6600 18236 -6572
rect 18476 -5748 19648 -5720
rect 18476 -6572 19564 -5748
rect 19628 -6572 19648 -5748
rect 18476 -6600 19648 -6572
rect 19888 -5748 21060 -5720
rect 19888 -6572 20976 -5748
rect 21040 -6572 21060 -5748
rect 19888 -6600 21060 -6572
rect 21300 -5748 22472 -5720
rect 21300 -6572 22388 -5748
rect 22452 -6572 22472 -5748
rect 21300 -6600 22472 -6572
rect 22712 -5748 23884 -5720
rect 22712 -6572 23800 -5748
rect 23864 -6572 23884 -5748
rect 22712 -6600 23884 -6572
rect -23884 -6868 -22712 -6840
rect -23884 -7692 -22796 -6868
rect -22732 -7692 -22712 -6868
rect -23884 -7720 -22712 -7692
rect -22472 -6868 -21300 -6840
rect -22472 -7692 -21384 -6868
rect -21320 -7692 -21300 -6868
rect -22472 -7720 -21300 -7692
rect -21060 -6868 -19888 -6840
rect -21060 -7692 -19972 -6868
rect -19908 -7692 -19888 -6868
rect -21060 -7720 -19888 -7692
rect -19648 -6868 -18476 -6840
rect -19648 -7692 -18560 -6868
rect -18496 -7692 -18476 -6868
rect -19648 -7720 -18476 -7692
rect -18236 -6868 -17064 -6840
rect -18236 -7692 -17148 -6868
rect -17084 -7692 -17064 -6868
rect -18236 -7720 -17064 -7692
rect -16824 -6868 -15652 -6840
rect -16824 -7692 -15736 -6868
rect -15672 -7692 -15652 -6868
rect -16824 -7720 -15652 -7692
rect -15412 -6868 -14240 -6840
rect -15412 -7692 -14324 -6868
rect -14260 -7692 -14240 -6868
rect -15412 -7720 -14240 -7692
rect -14000 -6868 -12828 -6840
rect -14000 -7692 -12912 -6868
rect -12848 -7692 -12828 -6868
rect -14000 -7720 -12828 -7692
rect -12588 -6868 -11416 -6840
rect -12588 -7692 -11500 -6868
rect -11436 -7692 -11416 -6868
rect -12588 -7720 -11416 -7692
rect -11176 -6868 -10004 -6840
rect -11176 -7692 -10088 -6868
rect -10024 -7692 -10004 -6868
rect -11176 -7720 -10004 -7692
rect -9764 -6868 -8592 -6840
rect -9764 -7692 -8676 -6868
rect -8612 -7692 -8592 -6868
rect -9764 -7720 -8592 -7692
rect -8352 -6868 -7180 -6840
rect -8352 -7692 -7264 -6868
rect -7200 -7692 -7180 -6868
rect -8352 -7720 -7180 -7692
rect -6940 -6868 -5768 -6840
rect -6940 -7692 -5852 -6868
rect -5788 -7692 -5768 -6868
rect -6940 -7720 -5768 -7692
rect -5528 -6868 -4356 -6840
rect -5528 -7692 -4440 -6868
rect -4376 -7692 -4356 -6868
rect -5528 -7720 -4356 -7692
rect -4116 -6868 -2944 -6840
rect -4116 -7692 -3028 -6868
rect -2964 -7692 -2944 -6868
rect -4116 -7720 -2944 -7692
rect -2704 -6868 -1532 -6840
rect -2704 -7692 -1616 -6868
rect -1552 -7692 -1532 -6868
rect -2704 -7720 -1532 -7692
rect -1292 -6868 -120 -6840
rect -1292 -7692 -204 -6868
rect -140 -7692 -120 -6868
rect -1292 -7720 -120 -7692
rect 120 -6868 1292 -6840
rect 120 -7692 1208 -6868
rect 1272 -7692 1292 -6868
rect 120 -7720 1292 -7692
rect 1532 -6868 2704 -6840
rect 1532 -7692 2620 -6868
rect 2684 -7692 2704 -6868
rect 1532 -7720 2704 -7692
rect 2944 -6868 4116 -6840
rect 2944 -7692 4032 -6868
rect 4096 -7692 4116 -6868
rect 2944 -7720 4116 -7692
rect 4356 -6868 5528 -6840
rect 4356 -7692 5444 -6868
rect 5508 -7692 5528 -6868
rect 4356 -7720 5528 -7692
rect 5768 -6868 6940 -6840
rect 5768 -7692 6856 -6868
rect 6920 -7692 6940 -6868
rect 5768 -7720 6940 -7692
rect 7180 -6868 8352 -6840
rect 7180 -7692 8268 -6868
rect 8332 -7692 8352 -6868
rect 7180 -7720 8352 -7692
rect 8592 -6868 9764 -6840
rect 8592 -7692 9680 -6868
rect 9744 -7692 9764 -6868
rect 8592 -7720 9764 -7692
rect 10004 -6868 11176 -6840
rect 10004 -7692 11092 -6868
rect 11156 -7692 11176 -6868
rect 10004 -7720 11176 -7692
rect 11416 -6868 12588 -6840
rect 11416 -7692 12504 -6868
rect 12568 -7692 12588 -6868
rect 11416 -7720 12588 -7692
rect 12828 -6868 14000 -6840
rect 12828 -7692 13916 -6868
rect 13980 -7692 14000 -6868
rect 12828 -7720 14000 -7692
rect 14240 -6868 15412 -6840
rect 14240 -7692 15328 -6868
rect 15392 -7692 15412 -6868
rect 14240 -7720 15412 -7692
rect 15652 -6868 16824 -6840
rect 15652 -7692 16740 -6868
rect 16804 -7692 16824 -6868
rect 15652 -7720 16824 -7692
rect 17064 -6868 18236 -6840
rect 17064 -7692 18152 -6868
rect 18216 -7692 18236 -6868
rect 17064 -7720 18236 -7692
rect 18476 -6868 19648 -6840
rect 18476 -7692 19564 -6868
rect 19628 -7692 19648 -6868
rect 18476 -7720 19648 -7692
rect 19888 -6868 21060 -6840
rect 19888 -7692 20976 -6868
rect 21040 -7692 21060 -6868
rect 19888 -7720 21060 -7692
rect 21300 -6868 22472 -6840
rect 21300 -7692 22388 -6868
rect 22452 -7692 22472 -6868
rect 21300 -7720 22472 -7692
rect 22712 -6868 23884 -6840
rect 22712 -7692 23800 -6868
rect 23864 -7692 23884 -6868
rect 22712 -7720 23884 -7692
rect -23884 -7988 -22712 -7960
rect -23884 -8812 -22796 -7988
rect -22732 -8812 -22712 -7988
rect -23884 -8840 -22712 -8812
rect -22472 -7988 -21300 -7960
rect -22472 -8812 -21384 -7988
rect -21320 -8812 -21300 -7988
rect -22472 -8840 -21300 -8812
rect -21060 -7988 -19888 -7960
rect -21060 -8812 -19972 -7988
rect -19908 -8812 -19888 -7988
rect -21060 -8840 -19888 -8812
rect -19648 -7988 -18476 -7960
rect -19648 -8812 -18560 -7988
rect -18496 -8812 -18476 -7988
rect -19648 -8840 -18476 -8812
rect -18236 -7988 -17064 -7960
rect -18236 -8812 -17148 -7988
rect -17084 -8812 -17064 -7988
rect -18236 -8840 -17064 -8812
rect -16824 -7988 -15652 -7960
rect -16824 -8812 -15736 -7988
rect -15672 -8812 -15652 -7988
rect -16824 -8840 -15652 -8812
rect -15412 -7988 -14240 -7960
rect -15412 -8812 -14324 -7988
rect -14260 -8812 -14240 -7988
rect -15412 -8840 -14240 -8812
rect -14000 -7988 -12828 -7960
rect -14000 -8812 -12912 -7988
rect -12848 -8812 -12828 -7988
rect -14000 -8840 -12828 -8812
rect -12588 -7988 -11416 -7960
rect -12588 -8812 -11500 -7988
rect -11436 -8812 -11416 -7988
rect -12588 -8840 -11416 -8812
rect -11176 -7988 -10004 -7960
rect -11176 -8812 -10088 -7988
rect -10024 -8812 -10004 -7988
rect -11176 -8840 -10004 -8812
rect -9764 -7988 -8592 -7960
rect -9764 -8812 -8676 -7988
rect -8612 -8812 -8592 -7988
rect -9764 -8840 -8592 -8812
rect -8352 -7988 -7180 -7960
rect -8352 -8812 -7264 -7988
rect -7200 -8812 -7180 -7988
rect -8352 -8840 -7180 -8812
rect -6940 -7988 -5768 -7960
rect -6940 -8812 -5852 -7988
rect -5788 -8812 -5768 -7988
rect -6940 -8840 -5768 -8812
rect -5528 -7988 -4356 -7960
rect -5528 -8812 -4440 -7988
rect -4376 -8812 -4356 -7988
rect -5528 -8840 -4356 -8812
rect -4116 -7988 -2944 -7960
rect -4116 -8812 -3028 -7988
rect -2964 -8812 -2944 -7988
rect -4116 -8840 -2944 -8812
rect -2704 -7988 -1532 -7960
rect -2704 -8812 -1616 -7988
rect -1552 -8812 -1532 -7988
rect -2704 -8840 -1532 -8812
rect -1292 -7988 -120 -7960
rect -1292 -8812 -204 -7988
rect -140 -8812 -120 -7988
rect -1292 -8840 -120 -8812
rect 120 -7988 1292 -7960
rect 120 -8812 1208 -7988
rect 1272 -8812 1292 -7988
rect 120 -8840 1292 -8812
rect 1532 -7988 2704 -7960
rect 1532 -8812 2620 -7988
rect 2684 -8812 2704 -7988
rect 1532 -8840 2704 -8812
rect 2944 -7988 4116 -7960
rect 2944 -8812 4032 -7988
rect 4096 -8812 4116 -7988
rect 2944 -8840 4116 -8812
rect 4356 -7988 5528 -7960
rect 4356 -8812 5444 -7988
rect 5508 -8812 5528 -7988
rect 4356 -8840 5528 -8812
rect 5768 -7988 6940 -7960
rect 5768 -8812 6856 -7988
rect 6920 -8812 6940 -7988
rect 5768 -8840 6940 -8812
rect 7180 -7988 8352 -7960
rect 7180 -8812 8268 -7988
rect 8332 -8812 8352 -7988
rect 7180 -8840 8352 -8812
rect 8592 -7988 9764 -7960
rect 8592 -8812 9680 -7988
rect 9744 -8812 9764 -7988
rect 8592 -8840 9764 -8812
rect 10004 -7988 11176 -7960
rect 10004 -8812 11092 -7988
rect 11156 -8812 11176 -7988
rect 10004 -8840 11176 -8812
rect 11416 -7988 12588 -7960
rect 11416 -8812 12504 -7988
rect 12568 -8812 12588 -7988
rect 11416 -8840 12588 -8812
rect 12828 -7988 14000 -7960
rect 12828 -8812 13916 -7988
rect 13980 -8812 14000 -7988
rect 12828 -8840 14000 -8812
rect 14240 -7988 15412 -7960
rect 14240 -8812 15328 -7988
rect 15392 -8812 15412 -7988
rect 14240 -8840 15412 -8812
rect 15652 -7988 16824 -7960
rect 15652 -8812 16740 -7988
rect 16804 -8812 16824 -7988
rect 15652 -8840 16824 -8812
rect 17064 -7988 18236 -7960
rect 17064 -8812 18152 -7988
rect 18216 -8812 18236 -7988
rect 17064 -8840 18236 -8812
rect 18476 -7988 19648 -7960
rect 18476 -8812 19564 -7988
rect 19628 -8812 19648 -7988
rect 18476 -8840 19648 -8812
rect 19888 -7988 21060 -7960
rect 19888 -8812 20976 -7988
rect 21040 -8812 21060 -7988
rect 19888 -8840 21060 -8812
rect 21300 -7988 22472 -7960
rect 21300 -8812 22388 -7988
rect 22452 -8812 22472 -7988
rect 21300 -8840 22472 -8812
rect 22712 -7988 23884 -7960
rect 22712 -8812 23800 -7988
rect 23864 -8812 23884 -7988
rect 22712 -8840 23884 -8812
rect -23884 -9108 -22712 -9080
rect -23884 -9932 -22796 -9108
rect -22732 -9932 -22712 -9108
rect -23884 -9960 -22712 -9932
rect -22472 -9108 -21300 -9080
rect -22472 -9932 -21384 -9108
rect -21320 -9932 -21300 -9108
rect -22472 -9960 -21300 -9932
rect -21060 -9108 -19888 -9080
rect -21060 -9932 -19972 -9108
rect -19908 -9932 -19888 -9108
rect -21060 -9960 -19888 -9932
rect -19648 -9108 -18476 -9080
rect -19648 -9932 -18560 -9108
rect -18496 -9932 -18476 -9108
rect -19648 -9960 -18476 -9932
rect -18236 -9108 -17064 -9080
rect -18236 -9932 -17148 -9108
rect -17084 -9932 -17064 -9108
rect -18236 -9960 -17064 -9932
rect -16824 -9108 -15652 -9080
rect -16824 -9932 -15736 -9108
rect -15672 -9932 -15652 -9108
rect -16824 -9960 -15652 -9932
rect -15412 -9108 -14240 -9080
rect -15412 -9932 -14324 -9108
rect -14260 -9932 -14240 -9108
rect -15412 -9960 -14240 -9932
rect -14000 -9108 -12828 -9080
rect -14000 -9932 -12912 -9108
rect -12848 -9932 -12828 -9108
rect -14000 -9960 -12828 -9932
rect -12588 -9108 -11416 -9080
rect -12588 -9932 -11500 -9108
rect -11436 -9932 -11416 -9108
rect -12588 -9960 -11416 -9932
rect -11176 -9108 -10004 -9080
rect -11176 -9932 -10088 -9108
rect -10024 -9932 -10004 -9108
rect -11176 -9960 -10004 -9932
rect -9764 -9108 -8592 -9080
rect -9764 -9932 -8676 -9108
rect -8612 -9932 -8592 -9108
rect -9764 -9960 -8592 -9932
rect -8352 -9108 -7180 -9080
rect -8352 -9932 -7264 -9108
rect -7200 -9932 -7180 -9108
rect -8352 -9960 -7180 -9932
rect -6940 -9108 -5768 -9080
rect -6940 -9932 -5852 -9108
rect -5788 -9932 -5768 -9108
rect -6940 -9960 -5768 -9932
rect -5528 -9108 -4356 -9080
rect -5528 -9932 -4440 -9108
rect -4376 -9932 -4356 -9108
rect -5528 -9960 -4356 -9932
rect -4116 -9108 -2944 -9080
rect -4116 -9932 -3028 -9108
rect -2964 -9932 -2944 -9108
rect -4116 -9960 -2944 -9932
rect -2704 -9108 -1532 -9080
rect -2704 -9932 -1616 -9108
rect -1552 -9932 -1532 -9108
rect -2704 -9960 -1532 -9932
rect -1292 -9108 -120 -9080
rect -1292 -9932 -204 -9108
rect -140 -9932 -120 -9108
rect -1292 -9960 -120 -9932
rect 120 -9108 1292 -9080
rect 120 -9932 1208 -9108
rect 1272 -9932 1292 -9108
rect 120 -9960 1292 -9932
rect 1532 -9108 2704 -9080
rect 1532 -9932 2620 -9108
rect 2684 -9932 2704 -9108
rect 1532 -9960 2704 -9932
rect 2944 -9108 4116 -9080
rect 2944 -9932 4032 -9108
rect 4096 -9932 4116 -9108
rect 2944 -9960 4116 -9932
rect 4356 -9108 5528 -9080
rect 4356 -9932 5444 -9108
rect 5508 -9932 5528 -9108
rect 4356 -9960 5528 -9932
rect 5768 -9108 6940 -9080
rect 5768 -9932 6856 -9108
rect 6920 -9932 6940 -9108
rect 5768 -9960 6940 -9932
rect 7180 -9108 8352 -9080
rect 7180 -9932 8268 -9108
rect 8332 -9932 8352 -9108
rect 7180 -9960 8352 -9932
rect 8592 -9108 9764 -9080
rect 8592 -9932 9680 -9108
rect 9744 -9932 9764 -9108
rect 8592 -9960 9764 -9932
rect 10004 -9108 11176 -9080
rect 10004 -9932 11092 -9108
rect 11156 -9932 11176 -9108
rect 10004 -9960 11176 -9932
rect 11416 -9108 12588 -9080
rect 11416 -9932 12504 -9108
rect 12568 -9932 12588 -9108
rect 11416 -9960 12588 -9932
rect 12828 -9108 14000 -9080
rect 12828 -9932 13916 -9108
rect 13980 -9932 14000 -9108
rect 12828 -9960 14000 -9932
rect 14240 -9108 15412 -9080
rect 14240 -9932 15328 -9108
rect 15392 -9932 15412 -9108
rect 14240 -9960 15412 -9932
rect 15652 -9108 16824 -9080
rect 15652 -9932 16740 -9108
rect 16804 -9932 16824 -9108
rect 15652 -9960 16824 -9932
rect 17064 -9108 18236 -9080
rect 17064 -9932 18152 -9108
rect 18216 -9932 18236 -9108
rect 17064 -9960 18236 -9932
rect 18476 -9108 19648 -9080
rect 18476 -9932 19564 -9108
rect 19628 -9932 19648 -9108
rect 18476 -9960 19648 -9932
rect 19888 -9108 21060 -9080
rect 19888 -9932 20976 -9108
rect 21040 -9932 21060 -9108
rect 19888 -9960 21060 -9932
rect 21300 -9108 22472 -9080
rect 21300 -9932 22388 -9108
rect 22452 -9932 22472 -9108
rect 21300 -9960 22472 -9932
rect 22712 -9108 23884 -9080
rect 22712 -9932 23800 -9108
rect 23864 -9932 23884 -9108
rect 22712 -9960 23884 -9932
rect -23884 -10228 -22712 -10200
rect -23884 -11052 -22796 -10228
rect -22732 -11052 -22712 -10228
rect -23884 -11080 -22712 -11052
rect -22472 -10228 -21300 -10200
rect -22472 -11052 -21384 -10228
rect -21320 -11052 -21300 -10228
rect -22472 -11080 -21300 -11052
rect -21060 -10228 -19888 -10200
rect -21060 -11052 -19972 -10228
rect -19908 -11052 -19888 -10228
rect -21060 -11080 -19888 -11052
rect -19648 -10228 -18476 -10200
rect -19648 -11052 -18560 -10228
rect -18496 -11052 -18476 -10228
rect -19648 -11080 -18476 -11052
rect -18236 -10228 -17064 -10200
rect -18236 -11052 -17148 -10228
rect -17084 -11052 -17064 -10228
rect -18236 -11080 -17064 -11052
rect -16824 -10228 -15652 -10200
rect -16824 -11052 -15736 -10228
rect -15672 -11052 -15652 -10228
rect -16824 -11080 -15652 -11052
rect -15412 -10228 -14240 -10200
rect -15412 -11052 -14324 -10228
rect -14260 -11052 -14240 -10228
rect -15412 -11080 -14240 -11052
rect -14000 -10228 -12828 -10200
rect -14000 -11052 -12912 -10228
rect -12848 -11052 -12828 -10228
rect -14000 -11080 -12828 -11052
rect -12588 -10228 -11416 -10200
rect -12588 -11052 -11500 -10228
rect -11436 -11052 -11416 -10228
rect -12588 -11080 -11416 -11052
rect -11176 -10228 -10004 -10200
rect -11176 -11052 -10088 -10228
rect -10024 -11052 -10004 -10228
rect -11176 -11080 -10004 -11052
rect -9764 -10228 -8592 -10200
rect -9764 -11052 -8676 -10228
rect -8612 -11052 -8592 -10228
rect -9764 -11080 -8592 -11052
rect -8352 -10228 -7180 -10200
rect -8352 -11052 -7264 -10228
rect -7200 -11052 -7180 -10228
rect -8352 -11080 -7180 -11052
rect -6940 -10228 -5768 -10200
rect -6940 -11052 -5852 -10228
rect -5788 -11052 -5768 -10228
rect -6940 -11080 -5768 -11052
rect -5528 -10228 -4356 -10200
rect -5528 -11052 -4440 -10228
rect -4376 -11052 -4356 -10228
rect -5528 -11080 -4356 -11052
rect -4116 -10228 -2944 -10200
rect -4116 -11052 -3028 -10228
rect -2964 -11052 -2944 -10228
rect -4116 -11080 -2944 -11052
rect -2704 -10228 -1532 -10200
rect -2704 -11052 -1616 -10228
rect -1552 -11052 -1532 -10228
rect -2704 -11080 -1532 -11052
rect -1292 -10228 -120 -10200
rect -1292 -11052 -204 -10228
rect -140 -11052 -120 -10228
rect -1292 -11080 -120 -11052
rect 120 -10228 1292 -10200
rect 120 -11052 1208 -10228
rect 1272 -11052 1292 -10228
rect 120 -11080 1292 -11052
rect 1532 -10228 2704 -10200
rect 1532 -11052 2620 -10228
rect 2684 -11052 2704 -10228
rect 1532 -11080 2704 -11052
rect 2944 -10228 4116 -10200
rect 2944 -11052 4032 -10228
rect 4096 -11052 4116 -10228
rect 2944 -11080 4116 -11052
rect 4356 -10228 5528 -10200
rect 4356 -11052 5444 -10228
rect 5508 -11052 5528 -10228
rect 4356 -11080 5528 -11052
rect 5768 -10228 6940 -10200
rect 5768 -11052 6856 -10228
rect 6920 -11052 6940 -10228
rect 5768 -11080 6940 -11052
rect 7180 -10228 8352 -10200
rect 7180 -11052 8268 -10228
rect 8332 -11052 8352 -10228
rect 7180 -11080 8352 -11052
rect 8592 -10228 9764 -10200
rect 8592 -11052 9680 -10228
rect 9744 -11052 9764 -10228
rect 8592 -11080 9764 -11052
rect 10004 -10228 11176 -10200
rect 10004 -11052 11092 -10228
rect 11156 -11052 11176 -10228
rect 10004 -11080 11176 -11052
rect 11416 -10228 12588 -10200
rect 11416 -11052 12504 -10228
rect 12568 -11052 12588 -10228
rect 11416 -11080 12588 -11052
rect 12828 -10228 14000 -10200
rect 12828 -11052 13916 -10228
rect 13980 -11052 14000 -10228
rect 12828 -11080 14000 -11052
rect 14240 -10228 15412 -10200
rect 14240 -11052 15328 -10228
rect 15392 -11052 15412 -10228
rect 14240 -11080 15412 -11052
rect 15652 -10228 16824 -10200
rect 15652 -11052 16740 -10228
rect 16804 -11052 16824 -10228
rect 15652 -11080 16824 -11052
rect 17064 -10228 18236 -10200
rect 17064 -11052 18152 -10228
rect 18216 -11052 18236 -10228
rect 17064 -11080 18236 -11052
rect 18476 -10228 19648 -10200
rect 18476 -11052 19564 -10228
rect 19628 -11052 19648 -10228
rect 18476 -11080 19648 -11052
rect 19888 -10228 21060 -10200
rect 19888 -11052 20976 -10228
rect 21040 -11052 21060 -10228
rect 19888 -11080 21060 -11052
rect 21300 -10228 22472 -10200
rect 21300 -11052 22388 -10228
rect 22452 -11052 22472 -10228
rect 21300 -11080 22472 -11052
rect 22712 -10228 23884 -10200
rect 22712 -11052 23800 -10228
rect 23864 -11052 23884 -10228
rect 22712 -11080 23884 -11052
rect -23884 -11348 -22712 -11320
rect -23884 -12172 -22796 -11348
rect -22732 -12172 -22712 -11348
rect -23884 -12200 -22712 -12172
rect -22472 -11348 -21300 -11320
rect -22472 -12172 -21384 -11348
rect -21320 -12172 -21300 -11348
rect -22472 -12200 -21300 -12172
rect -21060 -11348 -19888 -11320
rect -21060 -12172 -19972 -11348
rect -19908 -12172 -19888 -11348
rect -21060 -12200 -19888 -12172
rect -19648 -11348 -18476 -11320
rect -19648 -12172 -18560 -11348
rect -18496 -12172 -18476 -11348
rect -19648 -12200 -18476 -12172
rect -18236 -11348 -17064 -11320
rect -18236 -12172 -17148 -11348
rect -17084 -12172 -17064 -11348
rect -18236 -12200 -17064 -12172
rect -16824 -11348 -15652 -11320
rect -16824 -12172 -15736 -11348
rect -15672 -12172 -15652 -11348
rect -16824 -12200 -15652 -12172
rect -15412 -11348 -14240 -11320
rect -15412 -12172 -14324 -11348
rect -14260 -12172 -14240 -11348
rect -15412 -12200 -14240 -12172
rect -14000 -11348 -12828 -11320
rect -14000 -12172 -12912 -11348
rect -12848 -12172 -12828 -11348
rect -14000 -12200 -12828 -12172
rect -12588 -11348 -11416 -11320
rect -12588 -12172 -11500 -11348
rect -11436 -12172 -11416 -11348
rect -12588 -12200 -11416 -12172
rect -11176 -11348 -10004 -11320
rect -11176 -12172 -10088 -11348
rect -10024 -12172 -10004 -11348
rect -11176 -12200 -10004 -12172
rect -9764 -11348 -8592 -11320
rect -9764 -12172 -8676 -11348
rect -8612 -12172 -8592 -11348
rect -9764 -12200 -8592 -12172
rect -8352 -11348 -7180 -11320
rect -8352 -12172 -7264 -11348
rect -7200 -12172 -7180 -11348
rect -8352 -12200 -7180 -12172
rect -6940 -11348 -5768 -11320
rect -6940 -12172 -5852 -11348
rect -5788 -12172 -5768 -11348
rect -6940 -12200 -5768 -12172
rect -5528 -11348 -4356 -11320
rect -5528 -12172 -4440 -11348
rect -4376 -12172 -4356 -11348
rect -5528 -12200 -4356 -12172
rect -4116 -11348 -2944 -11320
rect -4116 -12172 -3028 -11348
rect -2964 -12172 -2944 -11348
rect -4116 -12200 -2944 -12172
rect -2704 -11348 -1532 -11320
rect -2704 -12172 -1616 -11348
rect -1552 -12172 -1532 -11348
rect -2704 -12200 -1532 -12172
rect -1292 -11348 -120 -11320
rect -1292 -12172 -204 -11348
rect -140 -12172 -120 -11348
rect -1292 -12200 -120 -12172
rect 120 -11348 1292 -11320
rect 120 -12172 1208 -11348
rect 1272 -12172 1292 -11348
rect 120 -12200 1292 -12172
rect 1532 -11348 2704 -11320
rect 1532 -12172 2620 -11348
rect 2684 -12172 2704 -11348
rect 1532 -12200 2704 -12172
rect 2944 -11348 4116 -11320
rect 2944 -12172 4032 -11348
rect 4096 -12172 4116 -11348
rect 2944 -12200 4116 -12172
rect 4356 -11348 5528 -11320
rect 4356 -12172 5444 -11348
rect 5508 -12172 5528 -11348
rect 4356 -12200 5528 -12172
rect 5768 -11348 6940 -11320
rect 5768 -12172 6856 -11348
rect 6920 -12172 6940 -11348
rect 5768 -12200 6940 -12172
rect 7180 -11348 8352 -11320
rect 7180 -12172 8268 -11348
rect 8332 -12172 8352 -11348
rect 7180 -12200 8352 -12172
rect 8592 -11348 9764 -11320
rect 8592 -12172 9680 -11348
rect 9744 -12172 9764 -11348
rect 8592 -12200 9764 -12172
rect 10004 -11348 11176 -11320
rect 10004 -12172 11092 -11348
rect 11156 -12172 11176 -11348
rect 10004 -12200 11176 -12172
rect 11416 -11348 12588 -11320
rect 11416 -12172 12504 -11348
rect 12568 -12172 12588 -11348
rect 11416 -12200 12588 -12172
rect 12828 -11348 14000 -11320
rect 12828 -12172 13916 -11348
rect 13980 -12172 14000 -11348
rect 12828 -12200 14000 -12172
rect 14240 -11348 15412 -11320
rect 14240 -12172 15328 -11348
rect 15392 -12172 15412 -11348
rect 14240 -12200 15412 -12172
rect 15652 -11348 16824 -11320
rect 15652 -12172 16740 -11348
rect 16804 -12172 16824 -11348
rect 15652 -12200 16824 -12172
rect 17064 -11348 18236 -11320
rect 17064 -12172 18152 -11348
rect 18216 -12172 18236 -11348
rect 17064 -12200 18236 -12172
rect 18476 -11348 19648 -11320
rect 18476 -12172 19564 -11348
rect 19628 -12172 19648 -11348
rect 18476 -12200 19648 -12172
rect 19888 -11348 21060 -11320
rect 19888 -12172 20976 -11348
rect 21040 -12172 21060 -11348
rect 19888 -12200 21060 -12172
rect 21300 -11348 22472 -11320
rect 21300 -12172 22388 -11348
rect 22452 -12172 22472 -11348
rect 21300 -12200 22472 -12172
rect 22712 -11348 23884 -11320
rect 22712 -12172 23800 -11348
rect 23864 -12172 23884 -11348
rect 22712 -12200 23884 -12172
rect -23884 -12468 -22712 -12440
rect -23884 -13292 -22796 -12468
rect -22732 -13292 -22712 -12468
rect -23884 -13320 -22712 -13292
rect -22472 -12468 -21300 -12440
rect -22472 -13292 -21384 -12468
rect -21320 -13292 -21300 -12468
rect -22472 -13320 -21300 -13292
rect -21060 -12468 -19888 -12440
rect -21060 -13292 -19972 -12468
rect -19908 -13292 -19888 -12468
rect -21060 -13320 -19888 -13292
rect -19648 -12468 -18476 -12440
rect -19648 -13292 -18560 -12468
rect -18496 -13292 -18476 -12468
rect -19648 -13320 -18476 -13292
rect -18236 -12468 -17064 -12440
rect -18236 -13292 -17148 -12468
rect -17084 -13292 -17064 -12468
rect -18236 -13320 -17064 -13292
rect -16824 -12468 -15652 -12440
rect -16824 -13292 -15736 -12468
rect -15672 -13292 -15652 -12468
rect -16824 -13320 -15652 -13292
rect -15412 -12468 -14240 -12440
rect -15412 -13292 -14324 -12468
rect -14260 -13292 -14240 -12468
rect -15412 -13320 -14240 -13292
rect -14000 -12468 -12828 -12440
rect -14000 -13292 -12912 -12468
rect -12848 -13292 -12828 -12468
rect -14000 -13320 -12828 -13292
rect -12588 -12468 -11416 -12440
rect -12588 -13292 -11500 -12468
rect -11436 -13292 -11416 -12468
rect -12588 -13320 -11416 -13292
rect -11176 -12468 -10004 -12440
rect -11176 -13292 -10088 -12468
rect -10024 -13292 -10004 -12468
rect -11176 -13320 -10004 -13292
rect -9764 -12468 -8592 -12440
rect -9764 -13292 -8676 -12468
rect -8612 -13292 -8592 -12468
rect -9764 -13320 -8592 -13292
rect -8352 -12468 -7180 -12440
rect -8352 -13292 -7264 -12468
rect -7200 -13292 -7180 -12468
rect -8352 -13320 -7180 -13292
rect -6940 -12468 -5768 -12440
rect -6940 -13292 -5852 -12468
rect -5788 -13292 -5768 -12468
rect -6940 -13320 -5768 -13292
rect -5528 -12468 -4356 -12440
rect -5528 -13292 -4440 -12468
rect -4376 -13292 -4356 -12468
rect -5528 -13320 -4356 -13292
rect -4116 -12468 -2944 -12440
rect -4116 -13292 -3028 -12468
rect -2964 -13292 -2944 -12468
rect -4116 -13320 -2944 -13292
rect -2704 -12468 -1532 -12440
rect -2704 -13292 -1616 -12468
rect -1552 -13292 -1532 -12468
rect -2704 -13320 -1532 -13292
rect -1292 -12468 -120 -12440
rect -1292 -13292 -204 -12468
rect -140 -13292 -120 -12468
rect -1292 -13320 -120 -13292
rect 120 -12468 1292 -12440
rect 120 -13292 1208 -12468
rect 1272 -13292 1292 -12468
rect 120 -13320 1292 -13292
rect 1532 -12468 2704 -12440
rect 1532 -13292 2620 -12468
rect 2684 -13292 2704 -12468
rect 1532 -13320 2704 -13292
rect 2944 -12468 4116 -12440
rect 2944 -13292 4032 -12468
rect 4096 -13292 4116 -12468
rect 2944 -13320 4116 -13292
rect 4356 -12468 5528 -12440
rect 4356 -13292 5444 -12468
rect 5508 -13292 5528 -12468
rect 4356 -13320 5528 -13292
rect 5768 -12468 6940 -12440
rect 5768 -13292 6856 -12468
rect 6920 -13292 6940 -12468
rect 5768 -13320 6940 -13292
rect 7180 -12468 8352 -12440
rect 7180 -13292 8268 -12468
rect 8332 -13292 8352 -12468
rect 7180 -13320 8352 -13292
rect 8592 -12468 9764 -12440
rect 8592 -13292 9680 -12468
rect 9744 -13292 9764 -12468
rect 8592 -13320 9764 -13292
rect 10004 -12468 11176 -12440
rect 10004 -13292 11092 -12468
rect 11156 -13292 11176 -12468
rect 10004 -13320 11176 -13292
rect 11416 -12468 12588 -12440
rect 11416 -13292 12504 -12468
rect 12568 -13292 12588 -12468
rect 11416 -13320 12588 -13292
rect 12828 -12468 14000 -12440
rect 12828 -13292 13916 -12468
rect 13980 -13292 14000 -12468
rect 12828 -13320 14000 -13292
rect 14240 -12468 15412 -12440
rect 14240 -13292 15328 -12468
rect 15392 -13292 15412 -12468
rect 14240 -13320 15412 -13292
rect 15652 -12468 16824 -12440
rect 15652 -13292 16740 -12468
rect 16804 -13292 16824 -12468
rect 15652 -13320 16824 -13292
rect 17064 -12468 18236 -12440
rect 17064 -13292 18152 -12468
rect 18216 -13292 18236 -12468
rect 17064 -13320 18236 -13292
rect 18476 -12468 19648 -12440
rect 18476 -13292 19564 -12468
rect 19628 -13292 19648 -12468
rect 18476 -13320 19648 -13292
rect 19888 -12468 21060 -12440
rect 19888 -13292 20976 -12468
rect 21040 -13292 21060 -12468
rect 19888 -13320 21060 -13292
rect 21300 -12468 22472 -12440
rect 21300 -13292 22388 -12468
rect 22452 -13292 22472 -12468
rect 21300 -13320 22472 -13292
rect 22712 -12468 23884 -12440
rect 22712 -13292 23800 -12468
rect 23864 -13292 23884 -12468
rect 22712 -13320 23884 -13292
rect -23884 -13588 -22712 -13560
rect -23884 -14412 -22796 -13588
rect -22732 -14412 -22712 -13588
rect -23884 -14440 -22712 -14412
rect -22472 -13588 -21300 -13560
rect -22472 -14412 -21384 -13588
rect -21320 -14412 -21300 -13588
rect -22472 -14440 -21300 -14412
rect -21060 -13588 -19888 -13560
rect -21060 -14412 -19972 -13588
rect -19908 -14412 -19888 -13588
rect -21060 -14440 -19888 -14412
rect -19648 -13588 -18476 -13560
rect -19648 -14412 -18560 -13588
rect -18496 -14412 -18476 -13588
rect -19648 -14440 -18476 -14412
rect -18236 -13588 -17064 -13560
rect -18236 -14412 -17148 -13588
rect -17084 -14412 -17064 -13588
rect -18236 -14440 -17064 -14412
rect -16824 -13588 -15652 -13560
rect -16824 -14412 -15736 -13588
rect -15672 -14412 -15652 -13588
rect -16824 -14440 -15652 -14412
rect -15412 -13588 -14240 -13560
rect -15412 -14412 -14324 -13588
rect -14260 -14412 -14240 -13588
rect -15412 -14440 -14240 -14412
rect -14000 -13588 -12828 -13560
rect -14000 -14412 -12912 -13588
rect -12848 -14412 -12828 -13588
rect -14000 -14440 -12828 -14412
rect -12588 -13588 -11416 -13560
rect -12588 -14412 -11500 -13588
rect -11436 -14412 -11416 -13588
rect -12588 -14440 -11416 -14412
rect -11176 -13588 -10004 -13560
rect -11176 -14412 -10088 -13588
rect -10024 -14412 -10004 -13588
rect -11176 -14440 -10004 -14412
rect -9764 -13588 -8592 -13560
rect -9764 -14412 -8676 -13588
rect -8612 -14412 -8592 -13588
rect -9764 -14440 -8592 -14412
rect -8352 -13588 -7180 -13560
rect -8352 -14412 -7264 -13588
rect -7200 -14412 -7180 -13588
rect -8352 -14440 -7180 -14412
rect -6940 -13588 -5768 -13560
rect -6940 -14412 -5852 -13588
rect -5788 -14412 -5768 -13588
rect -6940 -14440 -5768 -14412
rect -5528 -13588 -4356 -13560
rect -5528 -14412 -4440 -13588
rect -4376 -14412 -4356 -13588
rect -5528 -14440 -4356 -14412
rect -4116 -13588 -2944 -13560
rect -4116 -14412 -3028 -13588
rect -2964 -14412 -2944 -13588
rect -4116 -14440 -2944 -14412
rect -2704 -13588 -1532 -13560
rect -2704 -14412 -1616 -13588
rect -1552 -14412 -1532 -13588
rect -2704 -14440 -1532 -14412
rect -1292 -13588 -120 -13560
rect -1292 -14412 -204 -13588
rect -140 -14412 -120 -13588
rect -1292 -14440 -120 -14412
rect 120 -13588 1292 -13560
rect 120 -14412 1208 -13588
rect 1272 -14412 1292 -13588
rect 120 -14440 1292 -14412
rect 1532 -13588 2704 -13560
rect 1532 -14412 2620 -13588
rect 2684 -14412 2704 -13588
rect 1532 -14440 2704 -14412
rect 2944 -13588 4116 -13560
rect 2944 -14412 4032 -13588
rect 4096 -14412 4116 -13588
rect 2944 -14440 4116 -14412
rect 4356 -13588 5528 -13560
rect 4356 -14412 5444 -13588
rect 5508 -14412 5528 -13588
rect 4356 -14440 5528 -14412
rect 5768 -13588 6940 -13560
rect 5768 -14412 6856 -13588
rect 6920 -14412 6940 -13588
rect 5768 -14440 6940 -14412
rect 7180 -13588 8352 -13560
rect 7180 -14412 8268 -13588
rect 8332 -14412 8352 -13588
rect 7180 -14440 8352 -14412
rect 8592 -13588 9764 -13560
rect 8592 -14412 9680 -13588
rect 9744 -14412 9764 -13588
rect 8592 -14440 9764 -14412
rect 10004 -13588 11176 -13560
rect 10004 -14412 11092 -13588
rect 11156 -14412 11176 -13588
rect 10004 -14440 11176 -14412
rect 11416 -13588 12588 -13560
rect 11416 -14412 12504 -13588
rect 12568 -14412 12588 -13588
rect 11416 -14440 12588 -14412
rect 12828 -13588 14000 -13560
rect 12828 -14412 13916 -13588
rect 13980 -14412 14000 -13588
rect 12828 -14440 14000 -14412
rect 14240 -13588 15412 -13560
rect 14240 -14412 15328 -13588
rect 15392 -14412 15412 -13588
rect 14240 -14440 15412 -14412
rect 15652 -13588 16824 -13560
rect 15652 -14412 16740 -13588
rect 16804 -14412 16824 -13588
rect 15652 -14440 16824 -14412
rect 17064 -13588 18236 -13560
rect 17064 -14412 18152 -13588
rect 18216 -14412 18236 -13588
rect 17064 -14440 18236 -14412
rect 18476 -13588 19648 -13560
rect 18476 -14412 19564 -13588
rect 19628 -14412 19648 -13588
rect 18476 -14440 19648 -14412
rect 19888 -13588 21060 -13560
rect 19888 -14412 20976 -13588
rect 21040 -14412 21060 -13588
rect 19888 -14440 21060 -14412
rect 21300 -13588 22472 -13560
rect 21300 -14412 22388 -13588
rect 22452 -14412 22472 -13588
rect 21300 -14440 22472 -14412
rect 22712 -13588 23884 -13560
rect 22712 -14412 23800 -13588
rect 23864 -14412 23884 -13588
rect 22712 -14440 23884 -14412
rect -23884 -14708 -22712 -14680
rect -23884 -15532 -22796 -14708
rect -22732 -15532 -22712 -14708
rect -23884 -15560 -22712 -15532
rect -22472 -14708 -21300 -14680
rect -22472 -15532 -21384 -14708
rect -21320 -15532 -21300 -14708
rect -22472 -15560 -21300 -15532
rect -21060 -14708 -19888 -14680
rect -21060 -15532 -19972 -14708
rect -19908 -15532 -19888 -14708
rect -21060 -15560 -19888 -15532
rect -19648 -14708 -18476 -14680
rect -19648 -15532 -18560 -14708
rect -18496 -15532 -18476 -14708
rect -19648 -15560 -18476 -15532
rect -18236 -14708 -17064 -14680
rect -18236 -15532 -17148 -14708
rect -17084 -15532 -17064 -14708
rect -18236 -15560 -17064 -15532
rect -16824 -14708 -15652 -14680
rect -16824 -15532 -15736 -14708
rect -15672 -15532 -15652 -14708
rect -16824 -15560 -15652 -15532
rect -15412 -14708 -14240 -14680
rect -15412 -15532 -14324 -14708
rect -14260 -15532 -14240 -14708
rect -15412 -15560 -14240 -15532
rect -14000 -14708 -12828 -14680
rect -14000 -15532 -12912 -14708
rect -12848 -15532 -12828 -14708
rect -14000 -15560 -12828 -15532
rect -12588 -14708 -11416 -14680
rect -12588 -15532 -11500 -14708
rect -11436 -15532 -11416 -14708
rect -12588 -15560 -11416 -15532
rect -11176 -14708 -10004 -14680
rect -11176 -15532 -10088 -14708
rect -10024 -15532 -10004 -14708
rect -11176 -15560 -10004 -15532
rect -9764 -14708 -8592 -14680
rect -9764 -15532 -8676 -14708
rect -8612 -15532 -8592 -14708
rect -9764 -15560 -8592 -15532
rect -8352 -14708 -7180 -14680
rect -8352 -15532 -7264 -14708
rect -7200 -15532 -7180 -14708
rect -8352 -15560 -7180 -15532
rect -6940 -14708 -5768 -14680
rect -6940 -15532 -5852 -14708
rect -5788 -15532 -5768 -14708
rect -6940 -15560 -5768 -15532
rect -5528 -14708 -4356 -14680
rect -5528 -15532 -4440 -14708
rect -4376 -15532 -4356 -14708
rect -5528 -15560 -4356 -15532
rect -4116 -14708 -2944 -14680
rect -4116 -15532 -3028 -14708
rect -2964 -15532 -2944 -14708
rect -4116 -15560 -2944 -15532
rect -2704 -14708 -1532 -14680
rect -2704 -15532 -1616 -14708
rect -1552 -15532 -1532 -14708
rect -2704 -15560 -1532 -15532
rect -1292 -14708 -120 -14680
rect -1292 -15532 -204 -14708
rect -140 -15532 -120 -14708
rect -1292 -15560 -120 -15532
rect 120 -14708 1292 -14680
rect 120 -15532 1208 -14708
rect 1272 -15532 1292 -14708
rect 120 -15560 1292 -15532
rect 1532 -14708 2704 -14680
rect 1532 -15532 2620 -14708
rect 2684 -15532 2704 -14708
rect 1532 -15560 2704 -15532
rect 2944 -14708 4116 -14680
rect 2944 -15532 4032 -14708
rect 4096 -15532 4116 -14708
rect 2944 -15560 4116 -15532
rect 4356 -14708 5528 -14680
rect 4356 -15532 5444 -14708
rect 5508 -15532 5528 -14708
rect 4356 -15560 5528 -15532
rect 5768 -14708 6940 -14680
rect 5768 -15532 6856 -14708
rect 6920 -15532 6940 -14708
rect 5768 -15560 6940 -15532
rect 7180 -14708 8352 -14680
rect 7180 -15532 8268 -14708
rect 8332 -15532 8352 -14708
rect 7180 -15560 8352 -15532
rect 8592 -14708 9764 -14680
rect 8592 -15532 9680 -14708
rect 9744 -15532 9764 -14708
rect 8592 -15560 9764 -15532
rect 10004 -14708 11176 -14680
rect 10004 -15532 11092 -14708
rect 11156 -15532 11176 -14708
rect 10004 -15560 11176 -15532
rect 11416 -14708 12588 -14680
rect 11416 -15532 12504 -14708
rect 12568 -15532 12588 -14708
rect 11416 -15560 12588 -15532
rect 12828 -14708 14000 -14680
rect 12828 -15532 13916 -14708
rect 13980 -15532 14000 -14708
rect 12828 -15560 14000 -15532
rect 14240 -14708 15412 -14680
rect 14240 -15532 15328 -14708
rect 15392 -15532 15412 -14708
rect 14240 -15560 15412 -15532
rect 15652 -14708 16824 -14680
rect 15652 -15532 16740 -14708
rect 16804 -15532 16824 -14708
rect 15652 -15560 16824 -15532
rect 17064 -14708 18236 -14680
rect 17064 -15532 18152 -14708
rect 18216 -15532 18236 -14708
rect 17064 -15560 18236 -15532
rect 18476 -14708 19648 -14680
rect 18476 -15532 19564 -14708
rect 19628 -15532 19648 -14708
rect 18476 -15560 19648 -15532
rect 19888 -14708 21060 -14680
rect 19888 -15532 20976 -14708
rect 21040 -15532 21060 -14708
rect 19888 -15560 21060 -15532
rect 21300 -14708 22472 -14680
rect 21300 -15532 22388 -14708
rect 22452 -15532 22472 -14708
rect 21300 -15560 22472 -15532
rect 22712 -14708 23884 -14680
rect 22712 -15532 23800 -14708
rect 23864 -15532 23884 -14708
rect 22712 -15560 23884 -15532
rect -23884 -15828 -22712 -15800
rect -23884 -16652 -22796 -15828
rect -22732 -16652 -22712 -15828
rect -23884 -16680 -22712 -16652
rect -22472 -15828 -21300 -15800
rect -22472 -16652 -21384 -15828
rect -21320 -16652 -21300 -15828
rect -22472 -16680 -21300 -16652
rect -21060 -15828 -19888 -15800
rect -21060 -16652 -19972 -15828
rect -19908 -16652 -19888 -15828
rect -21060 -16680 -19888 -16652
rect -19648 -15828 -18476 -15800
rect -19648 -16652 -18560 -15828
rect -18496 -16652 -18476 -15828
rect -19648 -16680 -18476 -16652
rect -18236 -15828 -17064 -15800
rect -18236 -16652 -17148 -15828
rect -17084 -16652 -17064 -15828
rect -18236 -16680 -17064 -16652
rect -16824 -15828 -15652 -15800
rect -16824 -16652 -15736 -15828
rect -15672 -16652 -15652 -15828
rect -16824 -16680 -15652 -16652
rect -15412 -15828 -14240 -15800
rect -15412 -16652 -14324 -15828
rect -14260 -16652 -14240 -15828
rect -15412 -16680 -14240 -16652
rect -14000 -15828 -12828 -15800
rect -14000 -16652 -12912 -15828
rect -12848 -16652 -12828 -15828
rect -14000 -16680 -12828 -16652
rect -12588 -15828 -11416 -15800
rect -12588 -16652 -11500 -15828
rect -11436 -16652 -11416 -15828
rect -12588 -16680 -11416 -16652
rect -11176 -15828 -10004 -15800
rect -11176 -16652 -10088 -15828
rect -10024 -16652 -10004 -15828
rect -11176 -16680 -10004 -16652
rect -9764 -15828 -8592 -15800
rect -9764 -16652 -8676 -15828
rect -8612 -16652 -8592 -15828
rect -9764 -16680 -8592 -16652
rect -8352 -15828 -7180 -15800
rect -8352 -16652 -7264 -15828
rect -7200 -16652 -7180 -15828
rect -8352 -16680 -7180 -16652
rect -6940 -15828 -5768 -15800
rect -6940 -16652 -5852 -15828
rect -5788 -16652 -5768 -15828
rect -6940 -16680 -5768 -16652
rect -5528 -15828 -4356 -15800
rect -5528 -16652 -4440 -15828
rect -4376 -16652 -4356 -15828
rect -5528 -16680 -4356 -16652
rect -4116 -15828 -2944 -15800
rect -4116 -16652 -3028 -15828
rect -2964 -16652 -2944 -15828
rect -4116 -16680 -2944 -16652
rect -2704 -15828 -1532 -15800
rect -2704 -16652 -1616 -15828
rect -1552 -16652 -1532 -15828
rect -2704 -16680 -1532 -16652
rect -1292 -15828 -120 -15800
rect -1292 -16652 -204 -15828
rect -140 -16652 -120 -15828
rect -1292 -16680 -120 -16652
rect 120 -15828 1292 -15800
rect 120 -16652 1208 -15828
rect 1272 -16652 1292 -15828
rect 120 -16680 1292 -16652
rect 1532 -15828 2704 -15800
rect 1532 -16652 2620 -15828
rect 2684 -16652 2704 -15828
rect 1532 -16680 2704 -16652
rect 2944 -15828 4116 -15800
rect 2944 -16652 4032 -15828
rect 4096 -16652 4116 -15828
rect 2944 -16680 4116 -16652
rect 4356 -15828 5528 -15800
rect 4356 -16652 5444 -15828
rect 5508 -16652 5528 -15828
rect 4356 -16680 5528 -16652
rect 5768 -15828 6940 -15800
rect 5768 -16652 6856 -15828
rect 6920 -16652 6940 -15828
rect 5768 -16680 6940 -16652
rect 7180 -15828 8352 -15800
rect 7180 -16652 8268 -15828
rect 8332 -16652 8352 -15828
rect 7180 -16680 8352 -16652
rect 8592 -15828 9764 -15800
rect 8592 -16652 9680 -15828
rect 9744 -16652 9764 -15828
rect 8592 -16680 9764 -16652
rect 10004 -15828 11176 -15800
rect 10004 -16652 11092 -15828
rect 11156 -16652 11176 -15828
rect 10004 -16680 11176 -16652
rect 11416 -15828 12588 -15800
rect 11416 -16652 12504 -15828
rect 12568 -16652 12588 -15828
rect 11416 -16680 12588 -16652
rect 12828 -15828 14000 -15800
rect 12828 -16652 13916 -15828
rect 13980 -16652 14000 -15828
rect 12828 -16680 14000 -16652
rect 14240 -15828 15412 -15800
rect 14240 -16652 15328 -15828
rect 15392 -16652 15412 -15828
rect 14240 -16680 15412 -16652
rect 15652 -15828 16824 -15800
rect 15652 -16652 16740 -15828
rect 16804 -16652 16824 -15828
rect 15652 -16680 16824 -16652
rect 17064 -15828 18236 -15800
rect 17064 -16652 18152 -15828
rect 18216 -16652 18236 -15828
rect 17064 -16680 18236 -16652
rect 18476 -15828 19648 -15800
rect 18476 -16652 19564 -15828
rect 19628 -16652 19648 -15828
rect 18476 -16680 19648 -16652
rect 19888 -15828 21060 -15800
rect 19888 -16652 20976 -15828
rect 21040 -16652 21060 -15828
rect 19888 -16680 21060 -16652
rect 21300 -15828 22472 -15800
rect 21300 -16652 22388 -15828
rect 22452 -16652 22472 -15828
rect 21300 -16680 22472 -16652
rect 22712 -15828 23884 -15800
rect 22712 -16652 23800 -15828
rect 23864 -16652 23884 -15828
rect 22712 -16680 23884 -16652
rect -23884 -16948 -22712 -16920
rect -23884 -17772 -22796 -16948
rect -22732 -17772 -22712 -16948
rect -23884 -17800 -22712 -17772
rect -22472 -16948 -21300 -16920
rect -22472 -17772 -21384 -16948
rect -21320 -17772 -21300 -16948
rect -22472 -17800 -21300 -17772
rect -21060 -16948 -19888 -16920
rect -21060 -17772 -19972 -16948
rect -19908 -17772 -19888 -16948
rect -21060 -17800 -19888 -17772
rect -19648 -16948 -18476 -16920
rect -19648 -17772 -18560 -16948
rect -18496 -17772 -18476 -16948
rect -19648 -17800 -18476 -17772
rect -18236 -16948 -17064 -16920
rect -18236 -17772 -17148 -16948
rect -17084 -17772 -17064 -16948
rect -18236 -17800 -17064 -17772
rect -16824 -16948 -15652 -16920
rect -16824 -17772 -15736 -16948
rect -15672 -17772 -15652 -16948
rect -16824 -17800 -15652 -17772
rect -15412 -16948 -14240 -16920
rect -15412 -17772 -14324 -16948
rect -14260 -17772 -14240 -16948
rect -15412 -17800 -14240 -17772
rect -14000 -16948 -12828 -16920
rect -14000 -17772 -12912 -16948
rect -12848 -17772 -12828 -16948
rect -14000 -17800 -12828 -17772
rect -12588 -16948 -11416 -16920
rect -12588 -17772 -11500 -16948
rect -11436 -17772 -11416 -16948
rect -12588 -17800 -11416 -17772
rect -11176 -16948 -10004 -16920
rect -11176 -17772 -10088 -16948
rect -10024 -17772 -10004 -16948
rect -11176 -17800 -10004 -17772
rect -9764 -16948 -8592 -16920
rect -9764 -17772 -8676 -16948
rect -8612 -17772 -8592 -16948
rect -9764 -17800 -8592 -17772
rect -8352 -16948 -7180 -16920
rect -8352 -17772 -7264 -16948
rect -7200 -17772 -7180 -16948
rect -8352 -17800 -7180 -17772
rect -6940 -16948 -5768 -16920
rect -6940 -17772 -5852 -16948
rect -5788 -17772 -5768 -16948
rect -6940 -17800 -5768 -17772
rect -5528 -16948 -4356 -16920
rect -5528 -17772 -4440 -16948
rect -4376 -17772 -4356 -16948
rect -5528 -17800 -4356 -17772
rect -4116 -16948 -2944 -16920
rect -4116 -17772 -3028 -16948
rect -2964 -17772 -2944 -16948
rect -4116 -17800 -2944 -17772
rect -2704 -16948 -1532 -16920
rect -2704 -17772 -1616 -16948
rect -1552 -17772 -1532 -16948
rect -2704 -17800 -1532 -17772
rect -1292 -16948 -120 -16920
rect -1292 -17772 -204 -16948
rect -140 -17772 -120 -16948
rect -1292 -17800 -120 -17772
rect 120 -16948 1292 -16920
rect 120 -17772 1208 -16948
rect 1272 -17772 1292 -16948
rect 120 -17800 1292 -17772
rect 1532 -16948 2704 -16920
rect 1532 -17772 2620 -16948
rect 2684 -17772 2704 -16948
rect 1532 -17800 2704 -17772
rect 2944 -16948 4116 -16920
rect 2944 -17772 4032 -16948
rect 4096 -17772 4116 -16948
rect 2944 -17800 4116 -17772
rect 4356 -16948 5528 -16920
rect 4356 -17772 5444 -16948
rect 5508 -17772 5528 -16948
rect 4356 -17800 5528 -17772
rect 5768 -16948 6940 -16920
rect 5768 -17772 6856 -16948
rect 6920 -17772 6940 -16948
rect 5768 -17800 6940 -17772
rect 7180 -16948 8352 -16920
rect 7180 -17772 8268 -16948
rect 8332 -17772 8352 -16948
rect 7180 -17800 8352 -17772
rect 8592 -16948 9764 -16920
rect 8592 -17772 9680 -16948
rect 9744 -17772 9764 -16948
rect 8592 -17800 9764 -17772
rect 10004 -16948 11176 -16920
rect 10004 -17772 11092 -16948
rect 11156 -17772 11176 -16948
rect 10004 -17800 11176 -17772
rect 11416 -16948 12588 -16920
rect 11416 -17772 12504 -16948
rect 12568 -17772 12588 -16948
rect 11416 -17800 12588 -17772
rect 12828 -16948 14000 -16920
rect 12828 -17772 13916 -16948
rect 13980 -17772 14000 -16948
rect 12828 -17800 14000 -17772
rect 14240 -16948 15412 -16920
rect 14240 -17772 15328 -16948
rect 15392 -17772 15412 -16948
rect 14240 -17800 15412 -17772
rect 15652 -16948 16824 -16920
rect 15652 -17772 16740 -16948
rect 16804 -17772 16824 -16948
rect 15652 -17800 16824 -17772
rect 17064 -16948 18236 -16920
rect 17064 -17772 18152 -16948
rect 18216 -17772 18236 -16948
rect 17064 -17800 18236 -17772
rect 18476 -16948 19648 -16920
rect 18476 -17772 19564 -16948
rect 19628 -17772 19648 -16948
rect 18476 -17800 19648 -17772
rect 19888 -16948 21060 -16920
rect 19888 -17772 20976 -16948
rect 21040 -17772 21060 -16948
rect 19888 -17800 21060 -17772
rect 21300 -16948 22472 -16920
rect 21300 -17772 22388 -16948
rect 22452 -17772 22472 -16948
rect 21300 -17800 22472 -17772
rect 22712 -16948 23884 -16920
rect 22712 -17772 23800 -16948
rect 23864 -17772 23884 -16948
rect 22712 -17800 23884 -17772
rect -23884 -18068 -22712 -18040
rect -23884 -18892 -22796 -18068
rect -22732 -18892 -22712 -18068
rect -23884 -18920 -22712 -18892
rect -22472 -18068 -21300 -18040
rect -22472 -18892 -21384 -18068
rect -21320 -18892 -21300 -18068
rect -22472 -18920 -21300 -18892
rect -21060 -18068 -19888 -18040
rect -21060 -18892 -19972 -18068
rect -19908 -18892 -19888 -18068
rect -21060 -18920 -19888 -18892
rect -19648 -18068 -18476 -18040
rect -19648 -18892 -18560 -18068
rect -18496 -18892 -18476 -18068
rect -19648 -18920 -18476 -18892
rect -18236 -18068 -17064 -18040
rect -18236 -18892 -17148 -18068
rect -17084 -18892 -17064 -18068
rect -18236 -18920 -17064 -18892
rect -16824 -18068 -15652 -18040
rect -16824 -18892 -15736 -18068
rect -15672 -18892 -15652 -18068
rect -16824 -18920 -15652 -18892
rect -15412 -18068 -14240 -18040
rect -15412 -18892 -14324 -18068
rect -14260 -18892 -14240 -18068
rect -15412 -18920 -14240 -18892
rect -14000 -18068 -12828 -18040
rect -14000 -18892 -12912 -18068
rect -12848 -18892 -12828 -18068
rect -14000 -18920 -12828 -18892
rect -12588 -18068 -11416 -18040
rect -12588 -18892 -11500 -18068
rect -11436 -18892 -11416 -18068
rect -12588 -18920 -11416 -18892
rect -11176 -18068 -10004 -18040
rect -11176 -18892 -10088 -18068
rect -10024 -18892 -10004 -18068
rect -11176 -18920 -10004 -18892
rect -9764 -18068 -8592 -18040
rect -9764 -18892 -8676 -18068
rect -8612 -18892 -8592 -18068
rect -9764 -18920 -8592 -18892
rect -8352 -18068 -7180 -18040
rect -8352 -18892 -7264 -18068
rect -7200 -18892 -7180 -18068
rect -8352 -18920 -7180 -18892
rect -6940 -18068 -5768 -18040
rect -6940 -18892 -5852 -18068
rect -5788 -18892 -5768 -18068
rect -6940 -18920 -5768 -18892
rect -5528 -18068 -4356 -18040
rect -5528 -18892 -4440 -18068
rect -4376 -18892 -4356 -18068
rect -5528 -18920 -4356 -18892
rect -4116 -18068 -2944 -18040
rect -4116 -18892 -3028 -18068
rect -2964 -18892 -2944 -18068
rect -4116 -18920 -2944 -18892
rect -2704 -18068 -1532 -18040
rect -2704 -18892 -1616 -18068
rect -1552 -18892 -1532 -18068
rect -2704 -18920 -1532 -18892
rect -1292 -18068 -120 -18040
rect -1292 -18892 -204 -18068
rect -140 -18892 -120 -18068
rect -1292 -18920 -120 -18892
rect 120 -18068 1292 -18040
rect 120 -18892 1208 -18068
rect 1272 -18892 1292 -18068
rect 120 -18920 1292 -18892
rect 1532 -18068 2704 -18040
rect 1532 -18892 2620 -18068
rect 2684 -18892 2704 -18068
rect 1532 -18920 2704 -18892
rect 2944 -18068 4116 -18040
rect 2944 -18892 4032 -18068
rect 4096 -18892 4116 -18068
rect 2944 -18920 4116 -18892
rect 4356 -18068 5528 -18040
rect 4356 -18892 5444 -18068
rect 5508 -18892 5528 -18068
rect 4356 -18920 5528 -18892
rect 5768 -18068 6940 -18040
rect 5768 -18892 6856 -18068
rect 6920 -18892 6940 -18068
rect 5768 -18920 6940 -18892
rect 7180 -18068 8352 -18040
rect 7180 -18892 8268 -18068
rect 8332 -18892 8352 -18068
rect 7180 -18920 8352 -18892
rect 8592 -18068 9764 -18040
rect 8592 -18892 9680 -18068
rect 9744 -18892 9764 -18068
rect 8592 -18920 9764 -18892
rect 10004 -18068 11176 -18040
rect 10004 -18892 11092 -18068
rect 11156 -18892 11176 -18068
rect 10004 -18920 11176 -18892
rect 11416 -18068 12588 -18040
rect 11416 -18892 12504 -18068
rect 12568 -18892 12588 -18068
rect 11416 -18920 12588 -18892
rect 12828 -18068 14000 -18040
rect 12828 -18892 13916 -18068
rect 13980 -18892 14000 -18068
rect 12828 -18920 14000 -18892
rect 14240 -18068 15412 -18040
rect 14240 -18892 15328 -18068
rect 15392 -18892 15412 -18068
rect 14240 -18920 15412 -18892
rect 15652 -18068 16824 -18040
rect 15652 -18892 16740 -18068
rect 16804 -18892 16824 -18068
rect 15652 -18920 16824 -18892
rect 17064 -18068 18236 -18040
rect 17064 -18892 18152 -18068
rect 18216 -18892 18236 -18068
rect 17064 -18920 18236 -18892
rect 18476 -18068 19648 -18040
rect 18476 -18892 19564 -18068
rect 19628 -18892 19648 -18068
rect 18476 -18920 19648 -18892
rect 19888 -18068 21060 -18040
rect 19888 -18892 20976 -18068
rect 21040 -18892 21060 -18068
rect 19888 -18920 21060 -18892
rect 21300 -18068 22472 -18040
rect 21300 -18892 22388 -18068
rect 22452 -18892 22472 -18068
rect 21300 -18920 22472 -18892
rect 22712 -18068 23884 -18040
rect 22712 -18892 23800 -18068
rect 23864 -18892 23884 -18068
rect 22712 -18920 23884 -18892
<< via3 >>
rect -22796 18068 -22732 18892
rect -21384 18068 -21320 18892
rect -19972 18068 -19908 18892
rect -18560 18068 -18496 18892
rect -17148 18068 -17084 18892
rect -15736 18068 -15672 18892
rect -14324 18068 -14260 18892
rect -12912 18068 -12848 18892
rect -11500 18068 -11436 18892
rect -10088 18068 -10024 18892
rect -8676 18068 -8612 18892
rect -7264 18068 -7200 18892
rect -5852 18068 -5788 18892
rect -4440 18068 -4376 18892
rect -3028 18068 -2964 18892
rect -1616 18068 -1552 18892
rect -204 18068 -140 18892
rect 1208 18068 1272 18892
rect 2620 18068 2684 18892
rect 4032 18068 4096 18892
rect 5444 18068 5508 18892
rect 6856 18068 6920 18892
rect 8268 18068 8332 18892
rect 9680 18068 9744 18892
rect 11092 18068 11156 18892
rect 12504 18068 12568 18892
rect 13916 18068 13980 18892
rect 15328 18068 15392 18892
rect 16740 18068 16804 18892
rect 18152 18068 18216 18892
rect 19564 18068 19628 18892
rect 20976 18068 21040 18892
rect 22388 18068 22452 18892
rect 23800 18068 23864 18892
rect -22796 16948 -22732 17772
rect -21384 16948 -21320 17772
rect -19972 16948 -19908 17772
rect -18560 16948 -18496 17772
rect -17148 16948 -17084 17772
rect -15736 16948 -15672 17772
rect -14324 16948 -14260 17772
rect -12912 16948 -12848 17772
rect -11500 16948 -11436 17772
rect -10088 16948 -10024 17772
rect -8676 16948 -8612 17772
rect -7264 16948 -7200 17772
rect -5852 16948 -5788 17772
rect -4440 16948 -4376 17772
rect -3028 16948 -2964 17772
rect -1616 16948 -1552 17772
rect -204 16948 -140 17772
rect 1208 16948 1272 17772
rect 2620 16948 2684 17772
rect 4032 16948 4096 17772
rect 5444 16948 5508 17772
rect 6856 16948 6920 17772
rect 8268 16948 8332 17772
rect 9680 16948 9744 17772
rect 11092 16948 11156 17772
rect 12504 16948 12568 17772
rect 13916 16948 13980 17772
rect 15328 16948 15392 17772
rect 16740 16948 16804 17772
rect 18152 16948 18216 17772
rect 19564 16948 19628 17772
rect 20976 16948 21040 17772
rect 22388 16948 22452 17772
rect 23800 16948 23864 17772
rect -22796 15828 -22732 16652
rect -21384 15828 -21320 16652
rect -19972 15828 -19908 16652
rect -18560 15828 -18496 16652
rect -17148 15828 -17084 16652
rect -15736 15828 -15672 16652
rect -14324 15828 -14260 16652
rect -12912 15828 -12848 16652
rect -11500 15828 -11436 16652
rect -10088 15828 -10024 16652
rect -8676 15828 -8612 16652
rect -7264 15828 -7200 16652
rect -5852 15828 -5788 16652
rect -4440 15828 -4376 16652
rect -3028 15828 -2964 16652
rect -1616 15828 -1552 16652
rect -204 15828 -140 16652
rect 1208 15828 1272 16652
rect 2620 15828 2684 16652
rect 4032 15828 4096 16652
rect 5444 15828 5508 16652
rect 6856 15828 6920 16652
rect 8268 15828 8332 16652
rect 9680 15828 9744 16652
rect 11092 15828 11156 16652
rect 12504 15828 12568 16652
rect 13916 15828 13980 16652
rect 15328 15828 15392 16652
rect 16740 15828 16804 16652
rect 18152 15828 18216 16652
rect 19564 15828 19628 16652
rect 20976 15828 21040 16652
rect 22388 15828 22452 16652
rect 23800 15828 23864 16652
rect -22796 14708 -22732 15532
rect -21384 14708 -21320 15532
rect -19972 14708 -19908 15532
rect -18560 14708 -18496 15532
rect -17148 14708 -17084 15532
rect -15736 14708 -15672 15532
rect -14324 14708 -14260 15532
rect -12912 14708 -12848 15532
rect -11500 14708 -11436 15532
rect -10088 14708 -10024 15532
rect -8676 14708 -8612 15532
rect -7264 14708 -7200 15532
rect -5852 14708 -5788 15532
rect -4440 14708 -4376 15532
rect -3028 14708 -2964 15532
rect -1616 14708 -1552 15532
rect -204 14708 -140 15532
rect 1208 14708 1272 15532
rect 2620 14708 2684 15532
rect 4032 14708 4096 15532
rect 5444 14708 5508 15532
rect 6856 14708 6920 15532
rect 8268 14708 8332 15532
rect 9680 14708 9744 15532
rect 11092 14708 11156 15532
rect 12504 14708 12568 15532
rect 13916 14708 13980 15532
rect 15328 14708 15392 15532
rect 16740 14708 16804 15532
rect 18152 14708 18216 15532
rect 19564 14708 19628 15532
rect 20976 14708 21040 15532
rect 22388 14708 22452 15532
rect 23800 14708 23864 15532
rect -22796 13588 -22732 14412
rect -21384 13588 -21320 14412
rect -19972 13588 -19908 14412
rect -18560 13588 -18496 14412
rect -17148 13588 -17084 14412
rect -15736 13588 -15672 14412
rect -14324 13588 -14260 14412
rect -12912 13588 -12848 14412
rect -11500 13588 -11436 14412
rect -10088 13588 -10024 14412
rect -8676 13588 -8612 14412
rect -7264 13588 -7200 14412
rect -5852 13588 -5788 14412
rect -4440 13588 -4376 14412
rect -3028 13588 -2964 14412
rect -1616 13588 -1552 14412
rect -204 13588 -140 14412
rect 1208 13588 1272 14412
rect 2620 13588 2684 14412
rect 4032 13588 4096 14412
rect 5444 13588 5508 14412
rect 6856 13588 6920 14412
rect 8268 13588 8332 14412
rect 9680 13588 9744 14412
rect 11092 13588 11156 14412
rect 12504 13588 12568 14412
rect 13916 13588 13980 14412
rect 15328 13588 15392 14412
rect 16740 13588 16804 14412
rect 18152 13588 18216 14412
rect 19564 13588 19628 14412
rect 20976 13588 21040 14412
rect 22388 13588 22452 14412
rect 23800 13588 23864 14412
rect -22796 12468 -22732 13292
rect -21384 12468 -21320 13292
rect -19972 12468 -19908 13292
rect -18560 12468 -18496 13292
rect -17148 12468 -17084 13292
rect -15736 12468 -15672 13292
rect -14324 12468 -14260 13292
rect -12912 12468 -12848 13292
rect -11500 12468 -11436 13292
rect -10088 12468 -10024 13292
rect -8676 12468 -8612 13292
rect -7264 12468 -7200 13292
rect -5852 12468 -5788 13292
rect -4440 12468 -4376 13292
rect -3028 12468 -2964 13292
rect -1616 12468 -1552 13292
rect -204 12468 -140 13292
rect 1208 12468 1272 13292
rect 2620 12468 2684 13292
rect 4032 12468 4096 13292
rect 5444 12468 5508 13292
rect 6856 12468 6920 13292
rect 8268 12468 8332 13292
rect 9680 12468 9744 13292
rect 11092 12468 11156 13292
rect 12504 12468 12568 13292
rect 13916 12468 13980 13292
rect 15328 12468 15392 13292
rect 16740 12468 16804 13292
rect 18152 12468 18216 13292
rect 19564 12468 19628 13292
rect 20976 12468 21040 13292
rect 22388 12468 22452 13292
rect 23800 12468 23864 13292
rect -22796 11348 -22732 12172
rect -21384 11348 -21320 12172
rect -19972 11348 -19908 12172
rect -18560 11348 -18496 12172
rect -17148 11348 -17084 12172
rect -15736 11348 -15672 12172
rect -14324 11348 -14260 12172
rect -12912 11348 -12848 12172
rect -11500 11348 -11436 12172
rect -10088 11348 -10024 12172
rect -8676 11348 -8612 12172
rect -7264 11348 -7200 12172
rect -5852 11348 -5788 12172
rect -4440 11348 -4376 12172
rect -3028 11348 -2964 12172
rect -1616 11348 -1552 12172
rect -204 11348 -140 12172
rect 1208 11348 1272 12172
rect 2620 11348 2684 12172
rect 4032 11348 4096 12172
rect 5444 11348 5508 12172
rect 6856 11348 6920 12172
rect 8268 11348 8332 12172
rect 9680 11348 9744 12172
rect 11092 11348 11156 12172
rect 12504 11348 12568 12172
rect 13916 11348 13980 12172
rect 15328 11348 15392 12172
rect 16740 11348 16804 12172
rect 18152 11348 18216 12172
rect 19564 11348 19628 12172
rect 20976 11348 21040 12172
rect 22388 11348 22452 12172
rect 23800 11348 23864 12172
rect -22796 10228 -22732 11052
rect -21384 10228 -21320 11052
rect -19972 10228 -19908 11052
rect -18560 10228 -18496 11052
rect -17148 10228 -17084 11052
rect -15736 10228 -15672 11052
rect -14324 10228 -14260 11052
rect -12912 10228 -12848 11052
rect -11500 10228 -11436 11052
rect -10088 10228 -10024 11052
rect -8676 10228 -8612 11052
rect -7264 10228 -7200 11052
rect -5852 10228 -5788 11052
rect -4440 10228 -4376 11052
rect -3028 10228 -2964 11052
rect -1616 10228 -1552 11052
rect -204 10228 -140 11052
rect 1208 10228 1272 11052
rect 2620 10228 2684 11052
rect 4032 10228 4096 11052
rect 5444 10228 5508 11052
rect 6856 10228 6920 11052
rect 8268 10228 8332 11052
rect 9680 10228 9744 11052
rect 11092 10228 11156 11052
rect 12504 10228 12568 11052
rect 13916 10228 13980 11052
rect 15328 10228 15392 11052
rect 16740 10228 16804 11052
rect 18152 10228 18216 11052
rect 19564 10228 19628 11052
rect 20976 10228 21040 11052
rect 22388 10228 22452 11052
rect 23800 10228 23864 11052
rect -22796 9108 -22732 9932
rect -21384 9108 -21320 9932
rect -19972 9108 -19908 9932
rect -18560 9108 -18496 9932
rect -17148 9108 -17084 9932
rect -15736 9108 -15672 9932
rect -14324 9108 -14260 9932
rect -12912 9108 -12848 9932
rect -11500 9108 -11436 9932
rect -10088 9108 -10024 9932
rect -8676 9108 -8612 9932
rect -7264 9108 -7200 9932
rect -5852 9108 -5788 9932
rect -4440 9108 -4376 9932
rect -3028 9108 -2964 9932
rect -1616 9108 -1552 9932
rect -204 9108 -140 9932
rect 1208 9108 1272 9932
rect 2620 9108 2684 9932
rect 4032 9108 4096 9932
rect 5444 9108 5508 9932
rect 6856 9108 6920 9932
rect 8268 9108 8332 9932
rect 9680 9108 9744 9932
rect 11092 9108 11156 9932
rect 12504 9108 12568 9932
rect 13916 9108 13980 9932
rect 15328 9108 15392 9932
rect 16740 9108 16804 9932
rect 18152 9108 18216 9932
rect 19564 9108 19628 9932
rect 20976 9108 21040 9932
rect 22388 9108 22452 9932
rect 23800 9108 23864 9932
rect -22796 7988 -22732 8812
rect -21384 7988 -21320 8812
rect -19972 7988 -19908 8812
rect -18560 7988 -18496 8812
rect -17148 7988 -17084 8812
rect -15736 7988 -15672 8812
rect -14324 7988 -14260 8812
rect -12912 7988 -12848 8812
rect -11500 7988 -11436 8812
rect -10088 7988 -10024 8812
rect -8676 7988 -8612 8812
rect -7264 7988 -7200 8812
rect -5852 7988 -5788 8812
rect -4440 7988 -4376 8812
rect -3028 7988 -2964 8812
rect -1616 7988 -1552 8812
rect -204 7988 -140 8812
rect 1208 7988 1272 8812
rect 2620 7988 2684 8812
rect 4032 7988 4096 8812
rect 5444 7988 5508 8812
rect 6856 7988 6920 8812
rect 8268 7988 8332 8812
rect 9680 7988 9744 8812
rect 11092 7988 11156 8812
rect 12504 7988 12568 8812
rect 13916 7988 13980 8812
rect 15328 7988 15392 8812
rect 16740 7988 16804 8812
rect 18152 7988 18216 8812
rect 19564 7988 19628 8812
rect 20976 7988 21040 8812
rect 22388 7988 22452 8812
rect 23800 7988 23864 8812
rect -22796 6868 -22732 7692
rect -21384 6868 -21320 7692
rect -19972 6868 -19908 7692
rect -18560 6868 -18496 7692
rect -17148 6868 -17084 7692
rect -15736 6868 -15672 7692
rect -14324 6868 -14260 7692
rect -12912 6868 -12848 7692
rect -11500 6868 -11436 7692
rect -10088 6868 -10024 7692
rect -8676 6868 -8612 7692
rect -7264 6868 -7200 7692
rect -5852 6868 -5788 7692
rect -4440 6868 -4376 7692
rect -3028 6868 -2964 7692
rect -1616 6868 -1552 7692
rect -204 6868 -140 7692
rect 1208 6868 1272 7692
rect 2620 6868 2684 7692
rect 4032 6868 4096 7692
rect 5444 6868 5508 7692
rect 6856 6868 6920 7692
rect 8268 6868 8332 7692
rect 9680 6868 9744 7692
rect 11092 6868 11156 7692
rect 12504 6868 12568 7692
rect 13916 6868 13980 7692
rect 15328 6868 15392 7692
rect 16740 6868 16804 7692
rect 18152 6868 18216 7692
rect 19564 6868 19628 7692
rect 20976 6868 21040 7692
rect 22388 6868 22452 7692
rect 23800 6868 23864 7692
rect -22796 5748 -22732 6572
rect -21384 5748 -21320 6572
rect -19972 5748 -19908 6572
rect -18560 5748 -18496 6572
rect -17148 5748 -17084 6572
rect -15736 5748 -15672 6572
rect -14324 5748 -14260 6572
rect -12912 5748 -12848 6572
rect -11500 5748 -11436 6572
rect -10088 5748 -10024 6572
rect -8676 5748 -8612 6572
rect -7264 5748 -7200 6572
rect -5852 5748 -5788 6572
rect -4440 5748 -4376 6572
rect -3028 5748 -2964 6572
rect -1616 5748 -1552 6572
rect -204 5748 -140 6572
rect 1208 5748 1272 6572
rect 2620 5748 2684 6572
rect 4032 5748 4096 6572
rect 5444 5748 5508 6572
rect 6856 5748 6920 6572
rect 8268 5748 8332 6572
rect 9680 5748 9744 6572
rect 11092 5748 11156 6572
rect 12504 5748 12568 6572
rect 13916 5748 13980 6572
rect 15328 5748 15392 6572
rect 16740 5748 16804 6572
rect 18152 5748 18216 6572
rect 19564 5748 19628 6572
rect 20976 5748 21040 6572
rect 22388 5748 22452 6572
rect 23800 5748 23864 6572
rect -22796 4628 -22732 5452
rect -21384 4628 -21320 5452
rect -19972 4628 -19908 5452
rect -18560 4628 -18496 5452
rect -17148 4628 -17084 5452
rect -15736 4628 -15672 5452
rect -14324 4628 -14260 5452
rect -12912 4628 -12848 5452
rect -11500 4628 -11436 5452
rect -10088 4628 -10024 5452
rect -8676 4628 -8612 5452
rect -7264 4628 -7200 5452
rect -5852 4628 -5788 5452
rect -4440 4628 -4376 5452
rect -3028 4628 -2964 5452
rect -1616 4628 -1552 5452
rect -204 4628 -140 5452
rect 1208 4628 1272 5452
rect 2620 4628 2684 5452
rect 4032 4628 4096 5452
rect 5444 4628 5508 5452
rect 6856 4628 6920 5452
rect 8268 4628 8332 5452
rect 9680 4628 9744 5452
rect 11092 4628 11156 5452
rect 12504 4628 12568 5452
rect 13916 4628 13980 5452
rect 15328 4628 15392 5452
rect 16740 4628 16804 5452
rect 18152 4628 18216 5452
rect 19564 4628 19628 5452
rect 20976 4628 21040 5452
rect 22388 4628 22452 5452
rect 23800 4628 23864 5452
rect -22796 3508 -22732 4332
rect -21384 3508 -21320 4332
rect -19972 3508 -19908 4332
rect -18560 3508 -18496 4332
rect -17148 3508 -17084 4332
rect -15736 3508 -15672 4332
rect -14324 3508 -14260 4332
rect -12912 3508 -12848 4332
rect -11500 3508 -11436 4332
rect -10088 3508 -10024 4332
rect -8676 3508 -8612 4332
rect -7264 3508 -7200 4332
rect -5852 3508 -5788 4332
rect -4440 3508 -4376 4332
rect -3028 3508 -2964 4332
rect -1616 3508 -1552 4332
rect -204 3508 -140 4332
rect 1208 3508 1272 4332
rect 2620 3508 2684 4332
rect 4032 3508 4096 4332
rect 5444 3508 5508 4332
rect 6856 3508 6920 4332
rect 8268 3508 8332 4332
rect 9680 3508 9744 4332
rect 11092 3508 11156 4332
rect 12504 3508 12568 4332
rect 13916 3508 13980 4332
rect 15328 3508 15392 4332
rect 16740 3508 16804 4332
rect 18152 3508 18216 4332
rect 19564 3508 19628 4332
rect 20976 3508 21040 4332
rect 22388 3508 22452 4332
rect 23800 3508 23864 4332
rect -22796 2388 -22732 3212
rect -21384 2388 -21320 3212
rect -19972 2388 -19908 3212
rect -18560 2388 -18496 3212
rect -17148 2388 -17084 3212
rect -15736 2388 -15672 3212
rect -14324 2388 -14260 3212
rect -12912 2388 -12848 3212
rect -11500 2388 -11436 3212
rect -10088 2388 -10024 3212
rect -8676 2388 -8612 3212
rect -7264 2388 -7200 3212
rect -5852 2388 -5788 3212
rect -4440 2388 -4376 3212
rect -3028 2388 -2964 3212
rect -1616 2388 -1552 3212
rect -204 2388 -140 3212
rect 1208 2388 1272 3212
rect 2620 2388 2684 3212
rect 4032 2388 4096 3212
rect 5444 2388 5508 3212
rect 6856 2388 6920 3212
rect 8268 2388 8332 3212
rect 9680 2388 9744 3212
rect 11092 2388 11156 3212
rect 12504 2388 12568 3212
rect 13916 2388 13980 3212
rect 15328 2388 15392 3212
rect 16740 2388 16804 3212
rect 18152 2388 18216 3212
rect 19564 2388 19628 3212
rect 20976 2388 21040 3212
rect 22388 2388 22452 3212
rect 23800 2388 23864 3212
rect -22796 1268 -22732 2092
rect -21384 1268 -21320 2092
rect -19972 1268 -19908 2092
rect -18560 1268 -18496 2092
rect -17148 1268 -17084 2092
rect -15736 1268 -15672 2092
rect -14324 1268 -14260 2092
rect -12912 1268 -12848 2092
rect -11500 1268 -11436 2092
rect -10088 1268 -10024 2092
rect -8676 1268 -8612 2092
rect -7264 1268 -7200 2092
rect -5852 1268 -5788 2092
rect -4440 1268 -4376 2092
rect -3028 1268 -2964 2092
rect -1616 1268 -1552 2092
rect -204 1268 -140 2092
rect 1208 1268 1272 2092
rect 2620 1268 2684 2092
rect 4032 1268 4096 2092
rect 5444 1268 5508 2092
rect 6856 1268 6920 2092
rect 8268 1268 8332 2092
rect 9680 1268 9744 2092
rect 11092 1268 11156 2092
rect 12504 1268 12568 2092
rect 13916 1268 13980 2092
rect 15328 1268 15392 2092
rect 16740 1268 16804 2092
rect 18152 1268 18216 2092
rect 19564 1268 19628 2092
rect 20976 1268 21040 2092
rect 22388 1268 22452 2092
rect 23800 1268 23864 2092
rect -22796 148 -22732 972
rect -21384 148 -21320 972
rect -19972 148 -19908 972
rect -18560 148 -18496 972
rect -17148 148 -17084 972
rect -15736 148 -15672 972
rect -14324 148 -14260 972
rect -12912 148 -12848 972
rect -11500 148 -11436 972
rect -10088 148 -10024 972
rect -8676 148 -8612 972
rect -7264 148 -7200 972
rect -5852 148 -5788 972
rect -4440 148 -4376 972
rect -3028 148 -2964 972
rect -1616 148 -1552 972
rect -204 148 -140 972
rect 1208 148 1272 972
rect 2620 148 2684 972
rect 4032 148 4096 972
rect 5444 148 5508 972
rect 6856 148 6920 972
rect 8268 148 8332 972
rect 9680 148 9744 972
rect 11092 148 11156 972
rect 12504 148 12568 972
rect 13916 148 13980 972
rect 15328 148 15392 972
rect 16740 148 16804 972
rect 18152 148 18216 972
rect 19564 148 19628 972
rect 20976 148 21040 972
rect 22388 148 22452 972
rect 23800 148 23864 972
rect -22796 -972 -22732 -148
rect -21384 -972 -21320 -148
rect -19972 -972 -19908 -148
rect -18560 -972 -18496 -148
rect -17148 -972 -17084 -148
rect -15736 -972 -15672 -148
rect -14324 -972 -14260 -148
rect -12912 -972 -12848 -148
rect -11500 -972 -11436 -148
rect -10088 -972 -10024 -148
rect -8676 -972 -8612 -148
rect -7264 -972 -7200 -148
rect -5852 -972 -5788 -148
rect -4440 -972 -4376 -148
rect -3028 -972 -2964 -148
rect -1616 -972 -1552 -148
rect -204 -972 -140 -148
rect 1208 -972 1272 -148
rect 2620 -972 2684 -148
rect 4032 -972 4096 -148
rect 5444 -972 5508 -148
rect 6856 -972 6920 -148
rect 8268 -972 8332 -148
rect 9680 -972 9744 -148
rect 11092 -972 11156 -148
rect 12504 -972 12568 -148
rect 13916 -972 13980 -148
rect 15328 -972 15392 -148
rect 16740 -972 16804 -148
rect 18152 -972 18216 -148
rect 19564 -972 19628 -148
rect 20976 -972 21040 -148
rect 22388 -972 22452 -148
rect 23800 -972 23864 -148
rect -22796 -2092 -22732 -1268
rect -21384 -2092 -21320 -1268
rect -19972 -2092 -19908 -1268
rect -18560 -2092 -18496 -1268
rect -17148 -2092 -17084 -1268
rect -15736 -2092 -15672 -1268
rect -14324 -2092 -14260 -1268
rect -12912 -2092 -12848 -1268
rect -11500 -2092 -11436 -1268
rect -10088 -2092 -10024 -1268
rect -8676 -2092 -8612 -1268
rect -7264 -2092 -7200 -1268
rect -5852 -2092 -5788 -1268
rect -4440 -2092 -4376 -1268
rect -3028 -2092 -2964 -1268
rect -1616 -2092 -1552 -1268
rect -204 -2092 -140 -1268
rect 1208 -2092 1272 -1268
rect 2620 -2092 2684 -1268
rect 4032 -2092 4096 -1268
rect 5444 -2092 5508 -1268
rect 6856 -2092 6920 -1268
rect 8268 -2092 8332 -1268
rect 9680 -2092 9744 -1268
rect 11092 -2092 11156 -1268
rect 12504 -2092 12568 -1268
rect 13916 -2092 13980 -1268
rect 15328 -2092 15392 -1268
rect 16740 -2092 16804 -1268
rect 18152 -2092 18216 -1268
rect 19564 -2092 19628 -1268
rect 20976 -2092 21040 -1268
rect 22388 -2092 22452 -1268
rect 23800 -2092 23864 -1268
rect -22796 -3212 -22732 -2388
rect -21384 -3212 -21320 -2388
rect -19972 -3212 -19908 -2388
rect -18560 -3212 -18496 -2388
rect -17148 -3212 -17084 -2388
rect -15736 -3212 -15672 -2388
rect -14324 -3212 -14260 -2388
rect -12912 -3212 -12848 -2388
rect -11500 -3212 -11436 -2388
rect -10088 -3212 -10024 -2388
rect -8676 -3212 -8612 -2388
rect -7264 -3212 -7200 -2388
rect -5852 -3212 -5788 -2388
rect -4440 -3212 -4376 -2388
rect -3028 -3212 -2964 -2388
rect -1616 -3212 -1552 -2388
rect -204 -3212 -140 -2388
rect 1208 -3212 1272 -2388
rect 2620 -3212 2684 -2388
rect 4032 -3212 4096 -2388
rect 5444 -3212 5508 -2388
rect 6856 -3212 6920 -2388
rect 8268 -3212 8332 -2388
rect 9680 -3212 9744 -2388
rect 11092 -3212 11156 -2388
rect 12504 -3212 12568 -2388
rect 13916 -3212 13980 -2388
rect 15328 -3212 15392 -2388
rect 16740 -3212 16804 -2388
rect 18152 -3212 18216 -2388
rect 19564 -3212 19628 -2388
rect 20976 -3212 21040 -2388
rect 22388 -3212 22452 -2388
rect 23800 -3212 23864 -2388
rect -22796 -4332 -22732 -3508
rect -21384 -4332 -21320 -3508
rect -19972 -4332 -19908 -3508
rect -18560 -4332 -18496 -3508
rect -17148 -4332 -17084 -3508
rect -15736 -4332 -15672 -3508
rect -14324 -4332 -14260 -3508
rect -12912 -4332 -12848 -3508
rect -11500 -4332 -11436 -3508
rect -10088 -4332 -10024 -3508
rect -8676 -4332 -8612 -3508
rect -7264 -4332 -7200 -3508
rect -5852 -4332 -5788 -3508
rect -4440 -4332 -4376 -3508
rect -3028 -4332 -2964 -3508
rect -1616 -4332 -1552 -3508
rect -204 -4332 -140 -3508
rect 1208 -4332 1272 -3508
rect 2620 -4332 2684 -3508
rect 4032 -4332 4096 -3508
rect 5444 -4332 5508 -3508
rect 6856 -4332 6920 -3508
rect 8268 -4332 8332 -3508
rect 9680 -4332 9744 -3508
rect 11092 -4332 11156 -3508
rect 12504 -4332 12568 -3508
rect 13916 -4332 13980 -3508
rect 15328 -4332 15392 -3508
rect 16740 -4332 16804 -3508
rect 18152 -4332 18216 -3508
rect 19564 -4332 19628 -3508
rect 20976 -4332 21040 -3508
rect 22388 -4332 22452 -3508
rect 23800 -4332 23864 -3508
rect -22796 -5452 -22732 -4628
rect -21384 -5452 -21320 -4628
rect -19972 -5452 -19908 -4628
rect -18560 -5452 -18496 -4628
rect -17148 -5452 -17084 -4628
rect -15736 -5452 -15672 -4628
rect -14324 -5452 -14260 -4628
rect -12912 -5452 -12848 -4628
rect -11500 -5452 -11436 -4628
rect -10088 -5452 -10024 -4628
rect -8676 -5452 -8612 -4628
rect -7264 -5452 -7200 -4628
rect -5852 -5452 -5788 -4628
rect -4440 -5452 -4376 -4628
rect -3028 -5452 -2964 -4628
rect -1616 -5452 -1552 -4628
rect -204 -5452 -140 -4628
rect 1208 -5452 1272 -4628
rect 2620 -5452 2684 -4628
rect 4032 -5452 4096 -4628
rect 5444 -5452 5508 -4628
rect 6856 -5452 6920 -4628
rect 8268 -5452 8332 -4628
rect 9680 -5452 9744 -4628
rect 11092 -5452 11156 -4628
rect 12504 -5452 12568 -4628
rect 13916 -5452 13980 -4628
rect 15328 -5452 15392 -4628
rect 16740 -5452 16804 -4628
rect 18152 -5452 18216 -4628
rect 19564 -5452 19628 -4628
rect 20976 -5452 21040 -4628
rect 22388 -5452 22452 -4628
rect 23800 -5452 23864 -4628
rect -22796 -6572 -22732 -5748
rect -21384 -6572 -21320 -5748
rect -19972 -6572 -19908 -5748
rect -18560 -6572 -18496 -5748
rect -17148 -6572 -17084 -5748
rect -15736 -6572 -15672 -5748
rect -14324 -6572 -14260 -5748
rect -12912 -6572 -12848 -5748
rect -11500 -6572 -11436 -5748
rect -10088 -6572 -10024 -5748
rect -8676 -6572 -8612 -5748
rect -7264 -6572 -7200 -5748
rect -5852 -6572 -5788 -5748
rect -4440 -6572 -4376 -5748
rect -3028 -6572 -2964 -5748
rect -1616 -6572 -1552 -5748
rect -204 -6572 -140 -5748
rect 1208 -6572 1272 -5748
rect 2620 -6572 2684 -5748
rect 4032 -6572 4096 -5748
rect 5444 -6572 5508 -5748
rect 6856 -6572 6920 -5748
rect 8268 -6572 8332 -5748
rect 9680 -6572 9744 -5748
rect 11092 -6572 11156 -5748
rect 12504 -6572 12568 -5748
rect 13916 -6572 13980 -5748
rect 15328 -6572 15392 -5748
rect 16740 -6572 16804 -5748
rect 18152 -6572 18216 -5748
rect 19564 -6572 19628 -5748
rect 20976 -6572 21040 -5748
rect 22388 -6572 22452 -5748
rect 23800 -6572 23864 -5748
rect -22796 -7692 -22732 -6868
rect -21384 -7692 -21320 -6868
rect -19972 -7692 -19908 -6868
rect -18560 -7692 -18496 -6868
rect -17148 -7692 -17084 -6868
rect -15736 -7692 -15672 -6868
rect -14324 -7692 -14260 -6868
rect -12912 -7692 -12848 -6868
rect -11500 -7692 -11436 -6868
rect -10088 -7692 -10024 -6868
rect -8676 -7692 -8612 -6868
rect -7264 -7692 -7200 -6868
rect -5852 -7692 -5788 -6868
rect -4440 -7692 -4376 -6868
rect -3028 -7692 -2964 -6868
rect -1616 -7692 -1552 -6868
rect -204 -7692 -140 -6868
rect 1208 -7692 1272 -6868
rect 2620 -7692 2684 -6868
rect 4032 -7692 4096 -6868
rect 5444 -7692 5508 -6868
rect 6856 -7692 6920 -6868
rect 8268 -7692 8332 -6868
rect 9680 -7692 9744 -6868
rect 11092 -7692 11156 -6868
rect 12504 -7692 12568 -6868
rect 13916 -7692 13980 -6868
rect 15328 -7692 15392 -6868
rect 16740 -7692 16804 -6868
rect 18152 -7692 18216 -6868
rect 19564 -7692 19628 -6868
rect 20976 -7692 21040 -6868
rect 22388 -7692 22452 -6868
rect 23800 -7692 23864 -6868
rect -22796 -8812 -22732 -7988
rect -21384 -8812 -21320 -7988
rect -19972 -8812 -19908 -7988
rect -18560 -8812 -18496 -7988
rect -17148 -8812 -17084 -7988
rect -15736 -8812 -15672 -7988
rect -14324 -8812 -14260 -7988
rect -12912 -8812 -12848 -7988
rect -11500 -8812 -11436 -7988
rect -10088 -8812 -10024 -7988
rect -8676 -8812 -8612 -7988
rect -7264 -8812 -7200 -7988
rect -5852 -8812 -5788 -7988
rect -4440 -8812 -4376 -7988
rect -3028 -8812 -2964 -7988
rect -1616 -8812 -1552 -7988
rect -204 -8812 -140 -7988
rect 1208 -8812 1272 -7988
rect 2620 -8812 2684 -7988
rect 4032 -8812 4096 -7988
rect 5444 -8812 5508 -7988
rect 6856 -8812 6920 -7988
rect 8268 -8812 8332 -7988
rect 9680 -8812 9744 -7988
rect 11092 -8812 11156 -7988
rect 12504 -8812 12568 -7988
rect 13916 -8812 13980 -7988
rect 15328 -8812 15392 -7988
rect 16740 -8812 16804 -7988
rect 18152 -8812 18216 -7988
rect 19564 -8812 19628 -7988
rect 20976 -8812 21040 -7988
rect 22388 -8812 22452 -7988
rect 23800 -8812 23864 -7988
rect -22796 -9932 -22732 -9108
rect -21384 -9932 -21320 -9108
rect -19972 -9932 -19908 -9108
rect -18560 -9932 -18496 -9108
rect -17148 -9932 -17084 -9108
rect -15736 -9932 -15672 -9108
rect -14324 -9932 -14260 -9108
rect -12912 -9932 -12848 -9108
rect -11500 -9932 -11436 -9108
rect -10088 -9932 -10024 -9108
rect -8676 -9932 -8612 -9108
rect -7264 -9932 -7200 -9108
rect -5852 -9932 -5788 -9108
rect -4440 -9932 -4376 -9108
rect -3028 -9932 -2964 -9108
rect -1616 -9932 -1552 -9108
rect -204 -9932 -140 -9108
rect 1208 -9932 1272 -9108
rect 2620 -9932 2684 -9108
rect 4032 -9932 4096 -9108
rect 5444 -9932 5508 -9108
rect 6856 -9932 6920 -9108
rect 8268 -9932 8332 -9108
rect 9680 -9932 9744 -9108
rect 11092 -9932 11156 -9108
rect 12504 -9932 12568 -9108
rect 13916 -9932 13980 -9108
rect 15328 -9932 15392 -9108
rect 16740 -9932 16804 -9108
rect 18152 -9932 18216 -9108
rect 19564 -9932 19628 -9108
rect 20976 -9932 21040 -9108
rect 22388 -9932 22452 -9108
rect 23800 -9932 23864 -9108
rect -22796 -11052 -22732 -10228
rect -21384 -11052 -21320 -10228
rect -19972 -11052 -19908 -10228
rect -18560 -11052 -18496 -10228
rect -17148 -11052 -17084 -10228
rect -15736 -11052 -15672 -10228
rect -14324 -11052 -14260 -10228
rect -12912 -11052 -12848 -10228
rect -11500 -11052 -11436 -10228
rect -10088 -11052 -10024 -10228
rect -8676 -11052 -8612 -10228
rect -7264 -11052 -7200 -10228
rect -5852 -11052 -5788 -10228
rect -4440 -11052 -4376 -10228
rect -3028 -11052 -2964 -10228
rect -1616 -11052 -1552 -10228
rect -204 -11052 -140 -10228
rect 1208 -11052 1272 -10228
rect 2620 -11052 2684 -10228
rect 4032 -11052 4096 -10228
rect 5444 -11052 5508 -10228
rect 6856 -11052 6920 -10228
rect 8268 -11052 8332 -10228
rect 9680 -11052 9744 -10228
rect 11092 -11052 11156 -10228
rect 12504 -11052 12568 -10228
rect 13916 -11052 13980 -10228
rect 15328 -11052 15392 -10228
rect 16740 -11052 16804 -10228
rect 18152 -11052 18216 -10228
rect 19564 -11052 19628 -10228
rect 20976 -11052 21040 -10228
rect 22388 -11052 22452 -10228
rect 23800 -11052 23864 -10228
rect -22796 -12172 -22732 -11348
rect -21384 -12172 -21320 -11348
rect -19972 -12172 -19908 -11348
rect -18560 -12172 -18496 -11348
rect -17148 -12172 -17084 -11348
rect -15736 -12172 -15672 -11348
rect -14324 -12172 -14260 -11348
rect -12912 -12172 -12848 -11348
rect -11500 -12172 -11436 -11348
rect -10088 -12172 -10024 -11348
rect -8676 -12172 -8612 -11348
rect -7264 -12172 -7200 -11348
rect -5852 -12172 -5788 -11348
rect -4440 -12172 -4376 -11348
rect -3028 -12172 -2964 -11348
rect -1616 -12172 -1552 -11348
rect -204 -12172 -140 -11348
rect 1208 -12172 1272 -11348
rect 2620 -12172 2684 -11348
rect 4032 -12172 4096 -11348
rect 5444 -12172 5508 -11348
rect 6856 -12172 6920 -11348
rect 8268 -12172 8332 -11348
rect 9680 -12172 9744 -11348
rect 11092 -12172 11156 -11348
rect 12504 -12172 12568 -11348
rect 13916 -12172 13980 -11348
rect 15328 -12172 15392 -11348
rect 16740 -12172 16804 -11348
rect 18152 -12172 18216 -11348
rect 19564 -12172 19628 -11348
rect 20976 -12172 21040 -11348
rect 22388 -12172 22452 -11348
rect 23800 -12172 23864 -11348
rect -22796 -13292 -22732 -12468
rect -21384 -13292 -21320 -12468
rect -19972 -13292 -19908 -12468
rect -18560 -13292 -18496 -12468
rect -17148 -13292 -17084 -12468
rect -15736 -13292 -15672 -12468
rect -14324 -13292 -14260 -12468
rect -12912 -13292 -12848 -12468
rect -11500 -13292 -11436 -12468
rect -10088 -13292 -10024 -12468
rect -8676 -13292 -8612 -12468
rect -7264 -13292 -7200 -12468
rect -5852 -13292 -5788 -12468
rect -4440 -13292 -4376 -12468
rect -3028 -13292 -2964 -12468
rect -1616 -13292 -1552 -12468
rect -204 -13292 -140 -12468
rect 1208 -13292 1272 -12468
rect 2620 -13292 2684 -12468
rect 4032 -13292 4096 -12468
rect 5444 -13292 5508 -12468
rect 6856 -13292 6920 -12468
rect 8268 -13292 8332 -12468
rect 9680 -13292 9744 -12468
rect 11092 -13292 11156 -12468
rect 12504 -13292 12568 -12468
rect 13916 -13292 13980 -12468
rect 15328 -13292 15392 -12468
rect 16740 -13292 16804 -12468
rect 18152 -13292 18216 -12468
rect 19564 -13292 19628 -12468
rect 20976 -13292 21040 -12468
rect 22388 -13292 22452 -12468
rect 23800 -13292 23864 -12468
rect -22796 -14412 -22732 -13588
rect -21384 -14412 -21320 -13588
rect -19972 -14412 -19908 -13588
rect -18560 -14412 -18496 -13588
rect -17148 -14412 -17084 -13588
rect -15736 -14412 -15672 -13588
rect -14324 -14412 -14260 -13588
rect -12912 -14412 -12848 -13588
rect -11500 -14412 -11436 -13588
rect -10088 -14412 -10024 -13588
rect -8676 -14412 -8612 -13588
rect -7264 -14412 -7200 -13588
rect -5852 -14412 -5788 -13588
rect -4440 -14412 -4376 -13588
rect -3028 -14412 -2964 -13588
rect -1616 -14412 -1552 -13588
rect -204 -14412 -140 -13588
rect 1208 -14412 1272 -13588
rect 2620 -14412 2684 -13588
rect 4032 -14412 4096 -13588
rect 5444 -14412 5508 -13588
rect 6856 -14412 6920 -13588
rect 8268 -14412 8332 -13588
rect 9680 -14412 9744 -13588
rect 11092 -14412 11156 -13588
rect 12504 -14412 12568 -13588
rect 13916 -14412 13980 -13588
rect 15328 -14412 15392 -13588
rect 16740 -14412 16804 -13588
rect 18152 -14412 18216 -13588
rect 19564 -14412 19628 -13588
rect 20976 -14412 21040 -13588
rect 22388 -14412 22452 -13588
rect 23800 -14412 23864 -13588
rect -22796 -15532 -22732 -14708
rect -21384 -15532 -21320 -14708
rect -19972 -15532 -19908 -14708
rect -18560 -15532 -18496 -14708
rect -17148 -15532 -17084 -14708
rect -15736 -15532 -15672 -14708
rect -14324 -15532 -14260 -14708
rect -12912 -15532 -12848 -14708
rect -11500 -15532 -11436 -14708
rect -10088 -15532 -10024 -14708
rect -8676 -15532 -8612 -14708
rect -7264 -15532 -7200 -14708
rect -5852 -15532 -5788 -14708
rect -4440 -15532 -4376 -14708
rect -3028 -15532 -2964 -14708
rect -1616 -15532 -1552 -14708
rect -204 -15532 -140 -14708
rect 1208 -15532 1272 -14708
rect 2620 -15532 2684 -14708
rect 4032 -15532 4096 -14708
rect 5444 -15532 5508 -14708
rect 6856 -15532 6920 -14708
rect 8268 -15532 8332 -14708
rect 9680 -15532 9744 -14708
rect 11092 -15532 11156 -14708
rect 12504 -15532 12568 -14708
rect 13916 -15532 13980 -14708
rect 15328 -15532 15392 -14708
rect 16740 -15532 16804 -14708
rect 18152 -15532 18216 -14708
rect 19564 -15532 19628 -14708
rect 20976 -15532 21040 -14708
rect 22388 -15532 22452 -14708
rect 23800 -15532 23864 -14708
rect -22796 -16652 -22732 -15828
rect -21384 -16652 -21320 -15828
rect -19972 -16652 -19908 -15828
rect -18560 -16652 -18496 -15828
rect -17148 -16652 -17084 -15828
rect -15736 -16652 -15672 -15828
rect -14324 -16652 -14260 -15828
rect -12912 -16652 -12848 -15828
rect -11500 -16652 -11436 -15828
rect -10088 -16652 -10024 -15828
rect -8676 -16652 -8612 -15828
rect -7264 -16652 -7200 -15828
rect -5852 -16652 -5788 -15828
rect -4440 -16652 -4376 -15828
rect -3028 -16652 -2964 -15828
rect -1616 -16652 -1552 -15828
rect -204 -16652 -140 -15828
rect 1208 -16652 1272 -15828
rect 2620 -16652 2684 -15828
rect 4032 -16652 4096 -15828
rect 5444 -16652 5508 -15828
rect 6856 -16652 6920 -15828
rect 8268 -16652 8332 -15828
rect 9680 -16652 9744 -15828
rect 11092 -16652 11156 -15828
rect 12504 -16652 12568 -15828
rect 13916 -16652 13980 -15828
rect 15328 -16652 15392 -15828
rect 16740 -16652 16804 -15828
rect 18152 -16652 18216 -15828
rect 19564 -16652 19628 -15828
rect 20976 -16652 21040 -15828
rect 22388 -16652 22452 -15828
rect 23800 -16652 23864 -15828
rect -22796 -17772 -22732 -16948
rect -21384 -17772 -21320 -16948
rect -19972 -17772 -19908 -16948
rect -18560 -17772 -18496 -16948
rect -17148 -17772 -17084 -16948
rect -15736 -17772 -15672 -16948
rect -14324 -17772 -14260 -16948
rect -12912 -17772 -12848 -16948
rect -11500 -17772 -11436 -16948
rect -10088 -17772 -10024 -16948
rect -8676 -17772 -8612 -16948
rect -7264 -17772 -7200 -16948
rect -5852 -17772 -5788 -16948
rect -4440 -17772 -4376 -16948
rect -3028 -17772 -2964 -16948
rect -1616 -17772 -1552 -16948
rect -204 -17772 -140 -16948
rect 1208 -17772 1272 -16948
rect 2620 -17772 2684 -16948
rect 4032 -17772 4096 -16948
rect 5444 -17772 5508 -16948
rect 6856 -17772 6920 -16948
rect 8268 -17772 8332 -16948
rect 9680 -17772 9744 -16948
rect 11092 -17772 11156 -16948
rect 12504 -17772 12568 -16948
rect 13916 -17772 13980 -16948
rect 15328 -17772 15392 -16948
rect 16740 -17772 16804 -16948
rect 18152 -17772 18216 -16948
rect 19564 -17772 19628 -16948
rect 20976 -17772 21040 -16948
rect 22388 -17772 22452 -16948
rect 23800 -17772 23864 -16948
rect -22796 -18892 -22732 -18068
rect -21384 -18892 -21320 -18068
rect -19972 -18892 -19908 -18068
rect -18560 -18892 -18496 -18068
rect -17148 -18892 -17084 -18068
rect -15736 -18892 -15672 -18068
rect -14324 -18892 -14260 -18068
rect -12912 -18892 -12848 -18068
rect -11500 -18892 -11436 -18068
rect -10088 -18892 -10024 -18068
rect -8676 -18892 -8612 -18068
rect -7264 -18892 -7200 -18068
rect -5852 -18892 -5788 -18068
rect -4440 -18892 -4376 -18068
rect -3028 -18892 -2964 -18068
rect -1616 -18892 -1552 -18068
rect -204 -18892 -140 -18068
rect 1208 -18892 1272 -18068
rect 2620 -18892 2684 -18068
rect 4032 -18892 4096 -18068
rect 5444 -18892 5508 -18068
rect 6856 -18892 6920 -18068
rect 8268 -18892 8332 -18068
rect 9680 -18892 9744 -18068
rect 11092 -18892 11156 -18068
rect 12504 -18892 12568 -18068
rect 13916 -18892 13980 -18068
rect 15328 -18892 15392 -18068
rect 16740 -18892 16804 -18068
rect 18152 -18892 18216 -18068
rect 19564 -18892 19628 -18068
rect 20976 -18892 21040 -18068
rect 22388 -18892 22452 -18068
rect 23800 -18892 23864 -18068
<< mimcap >>
rect -23844 18840 -23044 18880
rect -23844 18120 -23804 18840
rect -23084 18120 -23044 18840
rect -23844 18080 -23044 18120
rect -22432 18840 -21632 18880
rect -22432 18120 -22392 18840
rect -21672 18120 -21632 18840
rect -22432 18080 -21632 18120
rect -21020 18840 -20220 18880
rect -21020 18120 -20980 18840
rect -20260 18120 -20220 18840
rect -21020 18080 -20220 18120
rect -19608 18840 -18808 18880
rect -19608 18120 -19568 18840
rect -18848 18120 -18808 18840
rect -19608 18080 -18808 18120
rect -18196 18840 -17396 18880
rect -18196 18120 -18156 18840
rect -17436 18120 -17396 18840
rect -18196 18080 -17396 18120
rect -16784 18840 -15984 18880
rect -16784 18120 -16744 18840
rect -16024 18120 -15984 18840
rect -16784 18080 -15984 18120
rect -15372 18840 -14572 18880
rect -15372 18120 -15332 18840
rect -14612 18120 -14572 18840
rect -15372 18080 -14572 18120
rect -13960 18840 -13160 18880
rect -13960 18120 -13920 18840
rect -13200 18120 -13160 18840
rect -13960 18080 -13160 18120
rect -12548 18840 -11748 18880
rect -12548 18120 -12508 18840
rect -11788 18120 -11748 18840
rect -12548 18080 -11748 18120
rect -11136 18840 -10336 18880
rect -11136 18120 -11096 18840
rect -10376 18120 -10336 18840
rect -11136 18080 -10336 18120
rect -9724 18840 -8924 18880
rect -9724 18120 -9684 18840
rect -8964 18120 -8924 18840
rect -9724 18080 -8924 18120
rect -8312 18840 -7512 18880
rect -8312 18120 -8272 18840
rect -7552 18120 -7512 18840
rect -8312 18080 -7512 18120
rect -6900 18840 -6100 18880
rect -6900 18120 -6860 18840
rect -6140 18120 -6100 18840
rect -6900 18080 -6100 18120
rect -5488 18840 -4688 18880
rect -5488 18120 -5448 18840
rect -4728 18120 -4688 18840
rect -5488 18080 -4688 18120
rect -4076 18840 -3276 18880
rect -4076 18120 -4036 18840
rect -3316 18120 -3276 18840
rect -4076 18080 -3276 18120
rect -2664 18840 -1864 18880
rect -2664 18120 -2624 18840
rect -1904 18120 -1864 18840
rect -2664 18080 -1864 18120
rect -1252 18840 -452 18880
rect -1252 18120 -1212 18840
rect -492 18120 -452 18840
rect -1252 18080 -452 18120
rect 160 18840 960 18880
rect 160 18120 200 18840
rect 920 18120 960 18840
rect 160 18080 960 18120
rect 1572 18840 2372 18880
rect 1572 18120 1612 18840
rect 2332 18120 2372 18840
rect 1572 18080 2372 18120
rect 2984 18840 3784 18880
rect 2984 18120 3024 18840
rect 3744 18120 3784 18840
rect 2984 18080 3784 18120
rect 4396 18840 5196 18880
rect 4396 18120 4436 18840
rect 5156 18120 5196 18840
rect 4396 18080 5196 18120
rect 5808 18840 6608 18880
rect 5808 18120 5848 18840
rect 6568 18120 6608 18840
rect 5808 18080 6608 18120
rect 7220 18840 8020 18880
rect 7220 18120 7260 18840
rect 7980 18120 8020 18840
rect 7220 18080 8020 18120
rect 8632 18840 9432 18880
rect 8632 18120 8672 18840
rect 9392 18120 9432 18840
rect 8632 18080 9432 18120
rect 10044 18840 10844 18880
rect 10044 18120 10084 18840
rect 10804 18120 10844 18840
rect 10044 18080 10844 18120
rect 11456 18840 12256 18880
rect 11456 18120 11496 18840
rect 12216 18120 12256 18840
rect 11456 18080 12256 18120
rect 12868 18840 13668 18880
rect 12868 18120 12908 18840
rect 13628 18120 13668 18840
rect 12868 18080 13668 18120
rect 14280 18840 15080 18880
rect 14280 18120 14320 18840
rect 15040 18120 15080 18840
rect 14280 18080 15080 18120
rect 15692 18840 16492 18880
rect 15692 18120 15732 18840
rect 16452 18120 16492 18840
rect 15692 18080 16492 18120
rect 17104 18840 17904 18880
rect 17104 18120 17144 18840
rect 17864 18120 17904 18840
rect 17104 18080 17904 18120
rect 18516 18840 19316 18880
rect 18516 18120 18556 18840
rect 19276 18120 19316 18840
rect 18516 18080 19316 18120
rect 19928 18840 20728 18880
rect 19928 18120 19968 18840
rect 20688 18120 20728 18840
rect 19928 18080 20728 18120
rect 21340 18840 22140 18880
rect 21340 18120 21380 18840
rect 22100 18120 22140 18840
rect 21340 18080 22140 18120
rect 22752 18840 23552 18880
rect 22752 18120 22792 18840
rect 23512 18120 23552 18840
rect 22752 18080 23552 18120
rect -23844 17720 -23044 17760
rect -23844 17000 -23804 17720
rect -23084 17000 -23044 17720
rect -23844 16960 -23044 17000
rect -22432 17720 -21632 17760
rect -22432 17000 -22392 17720
rect -21672 17000 -21632 17720
rect -22432 16960 -21632 17000
rect -21020 17720 -20220 17760
rect -21020 17000 -20980 17720
rect -20260 17000 -20220 17720
rect -21020 16960 -20220 17000
rect -19608 17720 -18808 17760
rect -19608 17000 -19568 17720
rect -18848 17000 -18808 17720
rect -19608 16960 -18808 17000
rect -18196 17720 -17396 17760
rect -18196 17000 -18156 17720
rect -17436 17000 -17396 17720
rect -18196 16960 -17396 17000
rect -16784 17720 -15984 17760
rect -16784 17000 -16744 17720
rect -16024 17000 -15984 17720
rect -16784 16960 -15984 17000
rect -15372 17720 -14572 17760
rect -15372 17000 -15332 17720
rect -14612 17000 -14572 17720
rect -15372 16960 -14572 17000
rect -13960 17720 -13160 17760
rect -13960 17000 -13920 17720
rect -13200 17000 -13160 17720
rect -13960 16960 -13160 17000
rect -12548 17720 -11748 17760
rect -12548 17000 -12508 17720
rect -11788 17000 -11748 17720
rect -12548 16960 -11748 17000
rect -11136 17720 -10336 17760
rect -11136 17000 -11096 17720
rect -10376 17000 -10336 17720
rect -11136 16960 -10336 17000
rect -9724 17720 -8924 17760
rect -9724 17000 -9684 17720
rect -8964 17000 -8924 17720
rect -9724 16960 -8924 17000
rect -8312 17720 -7512 17760
rect -8312 17000 -8272 17720
rect -7552 17000 -7512 17720
rect -8312 16960 -7512 17000
rect -6900 17720 -6100 17760
rect -6900 17000 -6860 17720
rect -6140 17000 -6100 17720
rect -6900 16960 -6100 17000
rect -5488 17720 -4688 17760
rect -5488 17000 -5448 17720
rect -4728 17000 -4688 17720
rect -5488 16960 -4688 17000
rect -4076 17720 -3276 17760
rect -4076 17000 -4036 17720
rect -3316 17000 -3276 17720
rect -4076 16960 -3276 17000
rect -2664 17720 -1864 17760
rect -2664 17000 -2624 17720
rect -1904 17000 -1864 17720
rect -2664 16960 -1864 17000
rect -1252 17720 -452 17760
rect -1252 17000 -1212 17720
rect -492 17000 -452 17720
rect -1252 16960 -452 17000
rect 160 17720 960 17760
rect 160 17000 200 17720
rect 920 17000 960 17720
rect 160 16960 960 17000
rect 1572 17720 2372 17760
rect 1572 17000 1612 17720
rect 2332 17000 2372 17720
rect 1572 16960 2372 17000
rect 2984 17720 3784 17760
rect 2984 17000 3024 17720
rect 3744 17000 3784 17720
rect 2984 16960 3784 17000
rect 4396 17720 5196 17760
rect 4396 17000 4436 17720
rect 5156 17000 5196 17720
rect 4396 16960 5196 17000
rect 5808 17720 6608 17760
rect 5808 17000 5848 17720
rect 6568 17000 6608 17720
rect 5808 16960 6608 17000
rect 7220 17720 8020 17760
rect 7220 17000 7260 17720
rect 7980 17000 8020 17720
rect 7220 16960 8020 17000
rect 8632 17720 9432 17760
rect 8632 17000 8672 17720
rect 9392 17000 9432 17720
rect 8632 16960 9432 17000
rect 10044 17720 10844 17760
rect 10044 17000 10084 17720
rect 10804 17000 10844 17720
rect 10044 16960 10844 17000
rect 11456 17720 12256 17760
rect 11456 17000 11496 17720
rect 12216 17000 12256 17720
rect 11456 16960 12256 17000
rect 12868 17720 13668 17760
rect 12868 17000 12908 17720
rect 13628 17000 13668 17720
rect 12868 16960 13668 17000
rect 14280 17720 15080 17760
rect 14280 17000 14320 17720
rect 15040 17000 15080 17720
rect 14280 16960 15080 17000
rect 15692 17720 16492 17760
rect 15692 17000 15732 17720
rect 16452 17000 16492 17720
rect 15692 16960 16492 17000
rect 17104 17720 17904 17760
rect 17104 17000 17144 17720
rect 17864 17000 17904 17720
rect 17104 16960 17904 17000
rect 18516 17720 19316 17760
rect 18516 17000 18556 17720
rect 19276 17000 19316 17720
rect 18516 16960 19316 17000
rect 19928 17720 20728 17760
rect 19928 17000 19968 17720
rect 20688 17000 20728 17720
rect 19928 16960 20728 17000
rect 21340 17720 22140 17760
rect 21340 17000 21380 17720
rect 22100 17000 22140 17720
rect 21340 16960 22140 17000
rect 22752 17720 23552 17760
rect 22752 17000 22792 17720
rect 23512 17000 23552 17720
rect 22752 16960 23552 17000
rect -23844 16600 -23044 16640
rect -23844 15880 -23804 16600
rect -23084 15880 -23044 16600
rect -23844 15840 -23044 15880
rect -22432 16600 -21632 16640
rect -22432 15880 -22392 16600
rect -21672 15880 -21632 16600
rect -22432 15840 -21632 15880
rect -21020 16600 -20220 16640
rect -21020 15880 -20980 16600
rect -20260 15880 -20220 16600
rect -21020 15840 -20220 15880
rect -19608 16600 -18808 16640
rect -19608 15880 -19568 16600
rect -18848 15880 -18808 16600
rect -19608 15840 -18808 15880
rect -18196 16600 -17396 16640
rect -18196 15880 -18156 16600
rect -17436 15880 -17396 16600
rect -18196 15840 -17396 15880
rect -16784 16600 -15984 16640
rect -16784 15880 -16744 16600
rect -16024 15880 -15984 16600
rect -16784 15840 -15984 15880
rect -15372 16600 -14572 16640
rect -15372 15880 -15332 16600
rect -14612 15880 -14572 16600
rect -15372 15840 -14572 15880
rect -13960 16600 -13160 16640
rect -13960 15880 -13920 16600
rect -13200 15880 -13160 16600
rect -13960 15840 -13160 15880
rect -12548 16600 -11748 16640
rect -12548 15880 -12508 16600
rect -11788 15880 -11748 16600
rect -12548 15840 -11748 15880
rect -11136 16600 -10336 16640
rect -11136 15880 -11096 16600
rect -10376 15880 -10336 16600
rect -11136 15840 -10336 15880
rect -9724 16600 -8924 16640
rect -9724 15880 -9684 16600
rect -8964 15880 -8924 16600
rect -9724 15840 -8924 15880
rect -8312 16600 -7512 16640
rect -8312 15880 -8272 16600
rect -7552 15880 -7512 16600
rect -8312 15840 -7512 15880
rect -6900 16600 -6100 16640
rect -6900 15880 -6860 16600
rect -6140 15880 -6100 16600
rect -6900 15840 -6100 15880
rect -5488 16600 -4688 16640
rect -5488 15880 -5448 16600
rect -4728 15880 -4688 16600
rect -5488 15840 -4688 15880
rect -4076 16600 -3276 16640
rect -4076 15880 -4036 16600
rect -3316 15880 -3276 16600
rect -4076 15840 -3276 15880
rect -2664 16600 -1864 16640
rect -2664 15880 -2624 16600
rect -1904 15880 -1864 16600
rect -2664 15840 -1864 15880
rect -1252 16600 -452 16640
rect -1252 15880 -1212 16600
rect -492 15880 -452 16600
rect -1252 15840 -452 15880
rect 160 16600 960 16640
rect 160 15880 200 16600
rect 920 15880 960 16600
rect 160 15840 960 15880
rect 1572 16600 2372 16640
rect 1572 15880 1612 16600
rect 2332 15880 2372 16600
rect 1572 15840 2372 15880
rect 2984 16600 3784 16640
rect 2984 15880 3024 16600
rect 3744 15880 3784 16600
rect 2984 15840 3784 15880
rect 4396 16600 5196 16640
rect 4396 15880 4436 16600
rect 5156 15880 5196 16600
rect 4396 15840 5196 15880
rect 5808 16600 6608 16640
rect 5808 15880 5848 16600
rect 6568 15880 6608 16600
rect 5808 15840 6608 15880
rect 7220 16600 8020 16640
rect 7220 15880 7260 16600
rect 7980 15880 8020 16600
rect 7220 15840 8020 15880
rect 8632 16600 9432 16640
rect 8632 15880 8672 16600
rect 9392 15880 9432 16600
rect 8632 15840 9432 15880
rect 10044 16600 10844 16640
rect 10044 15880 10084 16600
rect 10804 15880 10844 16600
rect 10044 15840 10844 15880
rect 11456 16600 12256 16640
rect 11456 15880 11496 16600
rect 12216 15880 12256 16600
rect 11456 15840 12256 15880
rect 12868 16600 13668 16640
rect 12868 15880 12908 16600
rect 13628 15880 13668 16600
rect 12868 15840 13668 15880
rect 14280 16600 15080 16640
rect 14280 15880 14320 16600
rect 15040 15880 15080 16600
rect 14280 15840 15080 15880
rect 15692 16600 16492 16640
rect 15692 15880 15732 16600
rect 16452 15880 16492 16600
rect 15692 15840 16492 15880
rect 17104 16600 17904 16640
rect 17104 15880 17144 16600
rect 17864 15880 17904 16600
rect 17104 15840 17904 15880
rect 18516 16600 19316 16640
rect 18516 15880 18556 16600
rect 19276 15880 19316 16600
rect 18516 15840 19316 15880
rect 19928 16600 20728 16640
rect 19928 15880 19968 16600
rect 20688 15880 20728 16600
rect 19928 15840 20728 15880
rect 21340 16600 22140 16640
rect 21340 15880 21380 16600
rect 22100 15880 22140 16600
rect 21340 15840 22140 15880
rect 22752 16600 23552 16640
rect 22752 15880 22792 16600
rect 23512 15880 23552 16600
rect 22752 15840 23552 15880
rect -23844 15480 -23044 15520
rect -23844 14760 -23804 15480
rect -23084 14760 -23044 15480
rect -23844 14720 -23044 14760
rect -22432 15480 -21632 15520
rect -22432 14760 -22392 15480
rect -21672 14760 -21632 15480
rect -22432 14720 -21632 14760
rect -21020 15480 -20220 15520
rect -21020 14760 -20980 15480
rect -20260 14760 -20220 15480
rect -21020 14720 -20220 14760
rect -19608 15480 -18808 15520
rect -19608 14760 -19568 15480
rect -18848 14760 -18808 15480
rect -19608 14720 -18808 14760
rect -18196 15480 -17396 15520
rect -18196 14760 -18156 15480
rect -17436 14760 -17396 15480
rect -18196 14720 -17396 14760
rect -16784 15480 -15984 15520
rect -16784 14760 -16744 15480
rect -16024 14760 -15984 15480
rect -16784 14720 -15984 14760
rect -15372 15480 -14572 15520
rect -15372 14760 -15332 15480
rect -14612 14760 -14572 15480
rect -15372 14720 -14572 14760
rect -13960 15480 -13160 15520
rect -13960 14760 -13920 15480
rect -13200 14760 -13160 15480
rect -13960 14720 -13160 14760
rect -12548 15480 -11748 15520
rect -12548 14760 -12508 15480
rect -11788 14760 -11748 15480
rect -12548 14720 -11748 14760
rect -11136 15480 -10336 15520
rect -11136 14760 -11096 15480
rect -10376 14760 -10336 15480
rect -11136 14720 -10336 14760
rect -9724 15480 -8924 15520
rect -9724 14760 -9684 15480
rect -8964 14760 -8924 15480
rect -9724 14720 -8924 14760
rect -8312 15480 -7512 15520
rect -8312 14760 -8272 15480
rect -7552 14760 -7512 15480
rect -8312 14720 -7512 14760
rect -6900 15480 -6100 15520
rect -6900 14760 -6860 15480
rect -6140 14760 -6100 15480
rect -6900 14720 -6100 14760
rect -5488 15480 -4688 15520
rect -5488 14760 -5448 15480
rect -4728 14760 -4688 15480
rect -5488 14720 -4688 14760
rect -4076 15480 -3276 15520
rect -4076 14760 -4036 15480
rect -3316 14760 -3276 15480
rect -4076 14720 -3276 14760
rect -2664 15480 -1864 15520
rect -2664 14760 -2624 15480
rect -1904 14760 -1864 15480
rect -2664 14720 -1864 14760
rect -1252 15480 -452 15520
rect -1252 14760 -1212 15480
rect -492 14760 -452 15480
rect -1252 14720 -452 14760
rect 160 15480 960 15520
rect 160 14760 200 15480
rect 920 14760 960 15480
rect 160 14720 960 14760
rect 1572 15480 2372 15520
rect 1572 14760 1612 15480
rect 2332 14760 2372 15480
rect 1572 14720 2372 14760
rect 2984 15480 3784 15520
rect 2984 14760 3024 15480
rect 3744 14760 3784 15480
rect 2984 14720 3784 14760
rect 4396 15480 5196 15520
rect 4396 14760 4436 15480
rect 5156 14760 5196 15480
rect 4396 14720 5196 14760
rect 5808 15480 6608 15520
rect 5808 14760 5848 15480
rect 6568 14760 6608 15480
rect 5808 14720 6608 14760
rect 7220 15480 8020 15520
rect 7220 14760 7260 15480
rect 7980 14760 8020 15480
rect 7220 14720 8020 14760
rect 8632 15480 9432 15520
rect 8632 14760 8672 15480
rect 9392 14760 9432 15480
rect 8632 14720 9432 14760
rect 10044 15480 10844 15520
rect 10044 14760 10084 15480
rect 10804 14760 10844 15480
rect 10044 14720 10844 14760
rect 11456 15480 12256 15520
rect 11456 14760 11496 15480
rect 12216 14760 12256 15480
rect 11456 14720 12256 14760
rect 12868 15480 13668 15520
rect 12868 14760 12908 15480
rect 13628 14760 13668 15480
rect 12868 14720 13668 14760
rect 14280 15480 15080 15520
rect 14280 14760 14320 15480
rect 15040 14760 15080 15480
rect 14280 14720 15080 14760
rect 15692 15480 16492 15520
rect 15692 14760 15732 15480
rect 16452 14760 16492 15480
rect 15692 14720 16492 14760
rect 17104 15480 17904 15520
rect 17104 14760 17144 15480
rect 17864 14760 17904 15480
rect 17104 14720 17904 14760
rect 18516 15480 19316 15520
rect 18516 14760 18556 15480
rect 19276 14760 19316 15480
rect 18516 14720 19316 14760
rect 19928 15480 20728 15520
rect 19928 14760 19968 15480
rect 20688 14760 20728 15480
rect 19928 14720 20728 14760
rect 21340 15480 22140 15520
rect 21340 14760 21380 15480
rect 22100 14760 22140 15480
rect 21340 14720 22140 14760
rect 22752 15480 23552 15520
rect 22752 14760 22792 15480
rect 23512 14760 23552 15480
rect 22752 14720 23552 14760
rect -23844 14360 -23044 14400
rect -23844 13640 -23804 14360
rect -23084 13640 -23044 14360
rect -23844 13600 -23044 13640
rect -22432 14360 -21632 14400
rect -22432 13640 -22392 14360
rect -21672 13640 -21632 14360
rect -22432 13600 -21632 13640
rect -21020 14360 -20220 14400
rect -21020 13640 -20980 14360
rect -20260 13640 -20220 14360
rect -21020 13600 -20220 13640
rect -19608 14360 -18808 14400
rect -19608 13640 -19568 14360
rect -18848 13640 -18808 14360
rect -19608 13600 -18808 13640
rect -18196 14360 -17396 14400
rect -18196 13640 -18156 14360
rect -17436 13640 -17396 14360
rect -18196 13600 -17396 13640
rect -16784 14360 -15984 14400
rect -16784 13640 -16744 14360
rect -16024 13640 -15984 14360
rect -16784 13600 -15984 13640
rect -15372 14360 -14572 14400
rect -15372 13640 -15332 14360
rect -14612 13640 -14572 14360
rect -15372 13600 -14572 13640
rect -13960 14360 -13160 14400
rect -13960 13640 -13920 14360
rect -13200 13640 -13160 14360
rect -13960 13600 -13160 13640
rect -12548 14360 -11748 14400
rect -12548 13640 -12508 14360
rect -11788 13640 -11748 14360
rect -12548 13600 -11748 13640
rect -11136 14360 -10336 14400
rect -11136 13640 -11096 14360
rect -10376 13640 -10336 14360
rect -11136 13600 -10336 13640
rect -9724 14360 -8924 14400
rect -9724 13640 -9684 14360
rect -8964 13640 -8924 14360
rect -9724 13600 -8924 13640
rect -8312 14360 -7512 14400
rect -8312 13640 -8272 14360
rect -7552 13640 -7512 14360
rect -8312 13600 -7512 13640
rect -6900 14360 -6100 14400
rect -6900 13640 -6860 14360
rect -6140 13640 -6100 14360
rect -6900 13600 -6100 13640
rect -5488 14360 -4688 14400
rect -5488 13640 -5448 14360
rect -4728 13640 -4688 14360
rect -5488 13600 -4688 13640
rect -4076 14360 -3276 14400
rect -4076 13640 -4036 14360
rect -3316 13640 -3276 14360
rect -4076 13600 -3276 13640
rect -2664 14360 -1864 14400
rect -2664 13640 -2624 14360
rect -1904 13640 -1864 14360
rect -2664 13600 -1864 13640
rect -1252 14360 -452 14400
rect -1252 13640 -1212 14360
rect -492 13640 -452 14360
rect -1252 13600 -452 13640
rect 160 14360 960 14400
rect 160 13640 200 14360
rect 920 13640 960 14360
rect 160 13600 960 13640
rect 1572 14360 2372 14400
rect 1572 13640 1612 14360
rect 2332 13640 2372 14360
rect 1572 13600 2372 13640
rect 2984 14360 3784 14400
rect 2984 13640 3024 14360
rect 3744 13640 3784 14360
rect 2984 13600 3784 13640
rect 4396 14360 5196 14400
rect 4396 13640 4436 14360
rect 5156 13640 5196 14360
rect 4396 13600 5196 13640
rect 5808 14360 6608 14400
rect 5808 13640 5848 14360
rect 6568 13640 6608 14360
rect 5808 13600 6608 13640
rect 7220 14360 8020 14400
rect 7220 13640 7260 14360
rect 7980 13640 8020 14360
rect 7220 13600 8020 13640
rect 8632 14360 9432 14400
rect 8632 13640 8672 14360
rect 9392 13640 9432 14360
rect 8632 13600 9432 13640
rect 10044 14360 10844 14400
rect 10044 13640 10084 14360
rect 10804 13640 10844 14360
rect 10044 13600 10844 13640
rect 11456 14360 12256 14400
rect 11456 13640 11496 14360
rect 12216 13640 12256 14360
rect 11456 13600 12256 13640
rect 12868 14360 13668 14400
rect 12868 13640 12908 14360
rect 13628 13640 13668 14360
rect 12868 13600 13668 13640
rect 14280 14360 15080 14400
rect 14280 13640 14320 14360
rect 15040 13640 15080 14360
rect 14280 13600 15080 13640
rect 15692 14360 16492 14400
rect 15692 13640 15732 14360
rect 16452 13640 16492 14360
rect 15692 13600 16492 13640
rect 17104 14360 17904 14400
rect 17104 13640 17144 14360
rect 17864 13640 17904 14360
rect 17104 13600 17904 13640
rect 18516 14360 19316 14400
rect 18516 13640 18556 14360
rect 19276 13640 19316 14360
rect 18516 13600 19316 13640
rect 19928 14360 20728 14400
rect 19928 13640 19968 14360
rect 20688 13640 20728 14360
rect 19928 13600 20728 13640
rect 21340 14360 22140 14400
rect 21340 13640 21380 14360
rect 22100 13640 22140 14360
rect 21340 13600 22140 13640
rect 22752 14360 23552 14400
rect 22752 13640 22792 14360
rect 23512 13640 23552 14360
rect 22752 13600 23552 13640
rect -23844 13240 -23044 13280
rect -23844 12520 -23804 13240
rect -23084 12520 -23044 13240
rect -23844 12480 -23044 12520
rect -22432 13240 -21632 13280
rect -22432 12520 -22392 13240
rect -21672 12520 -21632 13240
rect -22432 12480 -21632 12520
rect -21020 13240 -20220 13280
rect -21020 12520 -20980 13240
rect -20260 12520 -20220 13240
rect -21020 12480 -20220 12520
rect -19608 13240 -18808 13280
rect -19608 12520 -19568 13240
rect -18848 12520 -18808 13240
rect -19608 12480 -18808 12520
rect -18196 13240 -17396 13280
rect -18196 12520 -18156 13240
rect -17436 12520 -17396 13240
rect -18196 12480 -17396 12520
rect -16784 13240 -15984 13280
rect -16784 12520 -16744 13240
rect -16024 12520 -15984 13240
rect -16784 12480 -15984 12520
rect -15372 13240 -14572 13280
rect -15372 12520 -15332 13240
rect -14612 12520 -14572 13240
rect -15372 12480 -14572 12520
rect -13960 13240 -13160 13280
rect -13960 12520 -13920 13240
rect -13200 12520 -13160 13240
rect -13960 12480 -13160 12520
rect -12548 13240 -11748 13280
rect -12548 12520 -12508 13240
rect -11788 12520 -11748 13240
rect -12548 12480 -11748 12520
rect -11136 13240 -10336 13280
rect -11136 12520 -11096 13240
rect -10376 12520 -10336 13240
rect -11136 12480 -10336 12520
rect -9724 13240 -8924 13280
rect -9724 12520 -9684 13240
rect -8964 12520 -8924 13240
rect -9724 12480 -8924 12520
rect -8312 13240 -7512 13280
rect -8312 12520 -8272 13240
rect -7552 12520 -7512 13240
rect -8312 12480 -7512 12520
rect -6900 13240 -6100 13280
rect -6900 12520 -6860 13240
rect -6140 12520 -6100 13240
rect -6900 12480 -6100 12520
rect -5488 13240 -4688 13280
rect -5488 12520 -5448 13240
rect -4728 12520 -4688 13240
rect -5488 12480 -4688 12520
rect -4076 13240 -3276 13280
rect -4076 12520 -4036 13240
rect -3316 12520 -3276 13240
rect -4076 12480 -3276 12520
rect -2664 13240 -1864 13280
rect -2664 12520 -2624 13240
rect -1904 12520 -1864 13240
rect -2664 12480 -1864 12520
rect -1252 13240 -452 13280
rect -1252 12520 -1212 13240
rect -492 12520 -452 13240
rect -1252 12480 -452 12520
rect 160 13240 960 13280
rect 160 12520 200 13240
rect 920 12520 960 13240
rect 160 12480 960 12520
rect 1572 13240 2372 13280
rect 1572 12520 1612 13240
rect 2332 12520 2372 13240
rect 1572 12480 2372 12520
rect 2984 13240 3784 13280
rect 2984 12520 3024 13240
rect 3744 12520 3784 13240
rect 2984 12480 3784 12520
rect 4396 13240 5196 13280
rect 4396 12520 4436 13240
rect 5156 12520 5196 13240
rect 4396 12480 5196 12520
rect 5808 13240 6608 13280
rect 5808 12520 5848 13240
rect 6568 12520 6608 13240
rect 5808 12480 6608 12520
rect 7220 13240 8020 13280
rect 7220 12520 7260 13240
rect 7980 12520 8020 13240
rect 7220 12480 8020 12520
rect 8632 13240 9432 13280
rect 8632 12520 8672 13240
rect 9392 12520 9432 13240
rect 8632 12480 9432 12520
rect 10044 13240 10844 13280
rect 10044 12520 10084 13240
rect 10804 12520 10844 13240
rect 10044 12480 10844 12520
rect 11456 13240 12256 13280
rect 11456 12520 11496 13240
rect 12216 12520 12256 13240
rect 11456 12480 12256 12520
rect 12868 13240 13668 13280
rect 12868 12520 12908 13240
rect 13628 12520 13668 13240
rect 12868 12480 13668 12520
rect 14280 13240 15080 13280
rect 14280 12520 14320 13240
rect 15040 12520 15080 13240
rect 14280 12480 15080 12520
rect 15692 13240 16492 13280
rect 15692 12520 15732 13240
rect 16452 12520 16492 13240
rect 15692 12480 16492 12520
rect 17104 13240 17904 13280
rect 17104 12520 17144 13240
rect 17864 12520 17904 13240
rect 17104 12480 17904 12520
rect 18516 13240 19316 13280
rect 18516 12520 18556 13240
rect 19276 12520 19316 13240
rect 18516 12480 19316 12520
rect 19928 13240 20728 13280
rect 19928 12520 19968 13240
rect 20688 12520 20728 13240
rect 19928 12480 20728 12520
rect 21340 13240 22140 13280
rect 21340 12520 21380 13240
rect 22100 12520 22140 13240
rect 21340 12480 22140 12520
rect 22752 13240 23552 13280
rect 22752 12520 22792 13240
rect 23512 12520 23552 13240
rect 22752 12480 23552 12520
rect -23844 12120 -23044 12160
rect -23844 11400 -23804 12120
rect -23084 11400 -23044 12120
rect -23844 11360 -23044 11400
rect -22432 12120 -21632 12160
rect -22432 11400 -22392 12120
rect -21672 11400 -21632 12120
rect -22432 11360 -21632 11400
rect -21020 12120 -20220 12160
rect -21020 11400 -20980 12120
rect -20260 11400 -20220 12120
rect -21020 11360 -20220 11400
rect -19608 12120 -18808 12160
rect -19608 11400 -19568 12120
rect -18848 11400 -18808 12120
rect -19608 11360 -18808 11400
rect -18196 12120 -17396 12160
rect -18196 11400 -18156 12120
rect -17436 11400 -17396 12120
rect -18196 11360 -17396 11400
rect -16784 12120 -15984 12160
rect -16784 11400 -16744 12120
rect -16024 11400 -15984 12120
rect -16784 11360 -15984 11400
rect -15372 12120 -14572 12160
rect -15372 11400 -15332 12120
rect -14612 11400 -14572 12120
rect -15372 11360 -14572 11400
rect -13960 12120 -13160 12160
rect -13960 11400 -13920 12120
rect -13200 11400 -13160 12120
rect -13960 11360 -13160 11400
rect -12548 12120 -11748 12160
rect -12548 11400 -12508 12120
rect -11788 11400 -11748 12120
rect -12548 11360 -11748 11400
rect -11136 12120 -10336 12160
rect -11136 11400 -11096 12120
rect -10376 11400 -10336 12120
rect -11136 11360 -10336 11400
rect -9724 12120 -8924 12160
rect -9724 11400 -9684 12120
rect -8964 11400 -8924 12120
rect -9724 11360 -8924 11400
rect -8312 12120 -7512 12160
rect -8312 11400 -8272 12120
rect -7552 11400 -7512 12120
rect -8312 11360 -7512 11400
rect -6900 12120 -6100 12160
rect -6900 11400 -6860 12120
rect -6140 11400 -6100 12120
rect -6900 11360 -6100 11400
rect -5488 12120 -4688 12160
rect -5488 11400 -5448 12120
rect -4728 11400 -4688 12120
rect -5488 11360 -4688 11400
rect -4076 12120 -3276 12160
rect -4076 11400 -4036 12120
rect -3316 11400 -3276 12120
rect -4076 11360 -3276 11400
rect -2664 12120 -1864 12160
rect -2664 11400 -2624 12120
rect -1904 11400 -1864 12120
rect -2664 11360 -1864 11400
rect -1252 12120 -452 12160
rect -1252 11400 -1212 12120
rect -492 11400 -452 12120
rect -1252 11360 -452 11400
rect 160 12120 960 12160
rect 160 11400 200 12120
rect 920 11400 960 12120
rect 160 11360 960 11400
rect 1572 12120 2372 12160
rect 1572 11400 1612 12120
rect 2332 11400 2372 12120
rect 1572 11360 2372 11400
rect 2984 12120 3784 12160
rect 2984 11400 3024 12120
rect 3744 11400 3784 12120
rect 2984 11360 3784 11400
rect 4396 12120 5196 12160
rect 4396 11400 4436 12120
rect 5156 11400 5196 12120
rect 4396 11360 5196 11400
rect 5808 12120 6608 12160
rect 5808 11400 5848 12120
rect 6568 11400 6608 12120
rect 5808 11360 6608 11400
rect 7220 12120 8020 12160
rect 7220 11400 7260 12120
rect 7980 11400 8020 12120
rect 7220 11360 8020 11400
rect 8632 12120 9432 12160
rect 8632 11400 8672 12120
rect 9392 11400 9432 12120
rect 8632 11360 9432 11400
rect 10044 12120 10844 12160
rect 10044 11400 10084 12120
rect 10804 11400 10844 12120
rect 10044 11360 10844 11400
rect 11456 12120 12256 12160
rect 11456 11400 11496 12120
rect 12216 11400 12256 12120
rect 11456 11360 12256 11400
rect 12868 12120 13668 12160
rect 12868 11400 12908 12120
rect 13628 11400 13668 12120
rect 12868 11360 13668 11400
rect 14280 12120 15080 12160
rect 14280 11400 14320 12120
rect 15040 11400 15080 12120
rect 14280 11360 15080 11400
rect 15692 12120 16492 12160
rect 15692 11400 15732 12120
rect 16452 11400 16492 12120
rect 15692 11360 16492 11400
rect 17104 12120 17904 12160
rect 17104 11400 17144 12120
rect 17864 11400 17904 12120
rect 17104 11360 17904 11400
rect 18516 12120 19316 12160
rect 18516 11400 18556 12120
rect 19276 11400 19316 12120
rect 18516 11360 19316 11400
rect 19928 12120 20728 12160
rect 19928 11400 19968 12120
rect 20688 11400 20728 12120
rect 19928 11360 20728 11400
rect 21340 12120 22140 12160
rect 21340 11400 21380 12120
rect 22100 11400 22140 12120
rect 21340 11360 22140 11400
rect 22752 12120 23552 12160
rect 22752 11400 22792 12120
rect 23512 11400 23552 12120
rect 22752 11360 23552 11400
rect -23844 11000 -23044 11040
rect -23844 10280 -23804 11000
rect -23084 10280 -23044 11000
rect -23844 10240 -23044 10280
rect -22432 11000 -21632 11040
rect -22432 10280 -22392 11000
rect -21672 10280 -21632 11000
rect -22432 10240 -21632 10280
rect -21020 11000 -20220 11040
rect -21020 10280 -20980 11000
rect -20260 10280 -20220 11000
rect -21020 10240 -20220 10280
rect -19608 11000 -18808 11040
rect -19608 10280 -19568 11000
rect -18848 10280 -18808 11000
rect -19608 10240 -18808 10280
rect -18196 11000 -17396 11040
rect -18196 10280 -18156 11000
rect -17436 10280 -17396 11000
rect -18196 10240 -17396 10280
rect -16784 11000 -15984 11040
rect -16784 10280 -16744 11000
rect -16024 10280 -15984 11000
rect -16784 10240 -15984 10280
rect -15372 11000 -14572 11040
rect -15372 10280 -15332 11000
rect -14612 10280 -14572 11000
rect -15372 10240 -14572 10280
rect -13960 11000 -13160 11040
rect -13960 10280 -13920 11000
rect -13200 10280 -13160 11000
rect -13960 10240 -13160 10280
rect -12548 11000 -11748 11040
rect -12548 10280 -12508 11000
rect -11788 10280 -11748 11000
rect -12548 10240 -11748 10280
rect -11136 11000 -10336 11040
rect -11136 10280 -11096 11000
rect -10376 10280 -10336 11000
rect -11136 10240 -10336 10280
rect -9724 11000 -8924 11040
rect -9724 10280 -9684 11000
rect -8964 10280 -8924 11000
rect -9724 10240 -8924 10280
rect -8312 11000 -7512 11040
rect -8312 10280 -8272 11000
rect -7552 10280 -7512 11000
rect -8312 10240 -7512 10280
rect -6900 11000 -6100 11040
rect -6900 10280 -6860 11000
rect -6140 10280 -6100 11000
rect -6900 10240 -6100 10280
rect -5488 11000 -4688 11040
rect -5488 10280 -5448 11000
rect -4728 10280 -4688 11000
rect -5488 10240 -4688 10280
rect -4076 11000 -3276 11040
rect -4076 10280 -4036 11000
rect -3316 10280 -3276 11000
rect -4076 10240 -3276 10280
rect -2664 11000 -1864 11040
rect -2664 10280 -2624 11000
rect -1904 10280 -1864 11000
rect -2664 10240 -1864 10280
rect -1252 11000 -452 11040
rect -1252 10280 -1212 11000
rect -492 10280 -452 11000
rect -1252 10240 -452 10280
rect 160 11000 960 11040
rect 160 10280 200 11000
rect 920 10280 960 11000
rect 160 10240 960 10280
rect 1572 11000 2372 11040
rect 1572 10280 1612 11000
rect 2332 10280 2372 11000
rect 1572 10240 2372 10280
rect 2984 11000 3784 11040
rect 2984 10280 3024 11000
rect 3744 10280 3784 11000
rect 2984 10240 3784 10280
rect 4396 11000 5196 11040
rect 4396 10280 4436 11000
rect 5156 10280 5196 11000
rect 4396 10240 5196 10280
rect 5808 11000 6608 11040
rect 5808 10280 5848 11000
rect 6568 10280 6608 11000
rect 5808 10240 6608 10280
rect 7220 11000 8020 11040
rect 7220 10280 7260 11000
rect 7980 10280 8020 11000
rect 7220 10240 8020 10280
rect 8632 11000 9432 11040
rect 8632 10280 8672 11000
rect 9392 10280 9432 11000
rect 8632 10240 9432 10280
rect 10044 11000 10844 11040
rect 10044 10280 10084 11000
rect 10804 10280 10844 11000
rect 10044 10240 10844 10280
rect 11456 11000 12256 11040
rect 11456 10280 11496 11000
rect 12216 10280 12256 11000
rect 11456 10240 12256 10280
rect 12868 11000 13668 11040
rect 12868 10280 12908 11000
rect 13628 10280 13668 11000
rect 12868 10240 13668 10280
rect 14280 11000 15080 11040
rect 14280 10280 14320 11000
rect 15040 10280 15080 11000
rect 14280 10240 15080 10280
rect 15692 11000 16492 11040
rect 15692 10280 15732 11000
rect 16452 10280 16492 11000
rect 15692 10240 16492 10280
rect 17104 11000 17904 11040
rect 17104 10280 17144 11000
rect 17864 10280 17904 11000
rect 17104 10240 17904 10280
rect 18516 11000 19316 11040
rect 18516 10280 18556 11000
rect 19276 10280 19316 11000
rect 18516 10240 19316 10280
rect 19928 11000 20728 11040
rect 19928 10280 19968 11000
rect 20688 10280 20728 11000
rect 19928 10240 20728 10280
rect 21340 11000 22140 11040
rect 21340 10280 21380 11000
rect 22100 10280 22140 11000
rect 21340 10240 22140 10280
rect 22752 11000 23552 11040
rect 22752 10280 22792 11000
rect 23512 10280 23552 11000
rect 22752 10240 23552 10280
rect -23844 9880 -23044 9920
rect -23844 9160 -23804 9880
rect -23084 9160 -23044 9880
rect -23844 9120 -23044 9160
rect -22432 9880 -21632 9920
rect -22432 9160 -22392 9880
rect -21672 9160 -21632 9880
rect -22432 9120 -21632 9160
rect -21020 9880 -20220 9920
rect -21020 9160 -20980 9880
rect -20260 9160 -20220 9880
rect -21020 9120 -20220 9160
rect -19608 9880 -18808 9920
rect -19608 9160 -19568 9880
rect -18848 9160 -18808 9880
rect -19608 9120 -18808 9160
rect -18196 9880 -17396 9920
rect -18196 9160 -18156 9880
rect -17436 9160 -17396 9880
rect -18196 9120 -17396 9160
rect -16784 9880 -15984 9920
rect -16784 9160 -16744 9880
rect -16024 9160 -15984 9880
rect -16784 9120 -15984 9160
rect -15372 9880 -14572 9920
rect -15372 9160 -15332 9880
rect -14612 9160 -14572 9880
rect -15372 9120 -14572 9160
rect -13960 9880 -13160 9920
rect -13960 9160 -13920 9880
rect -13200 9160 -13160 9880
rect -13960 9120 -13160 9160
rect -12548 9880 -11748 9920
rect -12548 9160 -12508 9880
rect -11788 9160 -11748 9880
rect -12548 9120 -11748 9160
rect -11136 9880 -10336 9920
rect -11136 9160 -11096 9880
rect -10376 9160 -10336 9880
rect -11136 9120 -10336 9160
rect -9724 9880 -8924 9920
rect -9724 9160 -9684 9880
rect -8964 9160 -8924 9880
rect -9724 9120 -8924 9160
rect -8312 9880 -7512 9920
rect -8312 9160 -8272 9880
rect -7552 9160 -7512 9880
rect -8312 9120 -7512 9160
rect -6900 9880 -6100 9920
rect -6900 9160 -6860 9880
rect -6140 9160 -6100 9880
rect -6900 9120 -6100 9160
rect -5488 9880 -4688 9920
rect -5488 9160 -5448 9880
rect -4728 9160 -4688 9880
rect -5488 9120 -4688 9160
rect -4076 9880 -3276 9920
rect -4076 9160 -4036 9880
rect -3316 9160 -3276 9880
rect -4076 9120 -3276 9160
rect -2664 9880 -1864 9920
rect -2664 9160 -2624 9880
rect -1904 9160 -1864 9880
rect -2664 9120 -1864 9160
rect -1252 9880 -452 9920
rect -1252 9160 -1212 9880
rect -492 9160 -452 9880
rect -1252 9120 -452 9160
rect 160 9880 960 9920
rect 160 9160 200 9880
rect 920 9160 960 9880
rect 160 9120 960 9160
rect 1572 9880 2372 9920
rect 1572 9160 1612 9880
rect 2332 9160 2372 9880
rect 1572 9120 2372 9160
rect 2984 9880 3784 9920
rect 2984 9160 3024 9880
rect 3744 9160 3784 9880
rect 2984 9120 3784 9160
rect 4396 9880 5196 9920
rect 4396 9160 4436 9880
rect 5156 9160 5196 9880
rect 4396 9120 5196 9160
rect 5808 9880 6608 9920
rect 5808 9160 5848 9880
rect 6568 9160 6608 9880
rect 5808 9120 6608 9160
rect 7220 9880 8020 9920
rect 7220 9160 7260 9880
rect 7980 9160 8020 9880
rect 7220 9120 8020 9160
rect 8632 9880 9432 9920
rect 8632 9160 8672 9880
rect 9392 9160 9432 9880
rect 8632 9120 9432 9160
rect 10044 9880 10844 9920
rect 10044 9160 10084 9880
rect 10804 9160 10844 9880
rect 10044 9120 10844 9160
rect 11456 9880 12256 9920
rect 11456 9160 11496 9880
rect 12216 9160 12256 9880
rect 11456 9120 12256 9160
rect 12868 9880 13668 9920
rect 12868 9160 12908 9880
rect 13628 9160 13668 9880
rect 12868 9120 13668 9160
rect 14280 9880 15080 9920
rect 14280 9160 14320 9880
rect 15040 9160 15080 9880
rect 14280 9120 15080 9160
rect 15692 9880 16492 9920
rect 15692 9160 15732 9880
rect 16452 9160 16492 9880
rect 15692 9120 16492 9160
rect 17104 9880 17904 9920
rect 17104 9160 17144 9880
rect 17864 9160 17904 9880
rect 17104 9120 17904 9160
rect 18516 9880 19316 9920
rect 18516 9160 18556 9880
rect 19276 9160 19316 9880
rect 18516 9120 19316 9160
rect 19928 9880 20728 9920
rect 19928 9160 19968 9880
rect 20688 9160 20728 9880
rect 19928 9120 20728 9160
rect 21340 9880 22140 9920
rect 21340 9160 21380 9880
rect 22100 9160 22140 9880
rect 21340 9120 22140 9160
rect 22752 9880 23552 9920
rect 22752 9160 22792 9880
rect 23512 9160 23552 9880
rect 22752 9120 23552 9160
rect -23844 8760 -23044 8800
rect -23844 8040 -23804 8760
rect -23084 8040 -23044 8760
rect -23844 8000 -23044 8040
rect -22432 8760 -21632 8800
rect -22432 8040 -22392 8760
rect -21672 8040 -21632 8760
rect -22432 8000 -21632 8040
rect -21020 8760 -20220 8800
rect -21020 8040 -20980 8760
rect -20260 8040 -20220 8760
rect -21020 8000 -20220 8040
rect -19608 8760 -18808 8800
rect -19608 8040 -19568 8760
rect -18848 8040 -18808 8760
rect -19608 8000 -18808 8040
rect -18196 8760 -17396 8800
rect -18196 8040 -18156 8760
rect -17436 8040 -17396 8760
rect -18196 8000 -17396 8040
rect -16784 8760 -15984 8800
rect -16784 8040 -16744 8760
rect -16024 8040 -15984 8760
rect -16784 8000 -15984 8040
rect -15372 8760 -14572 8800
rect -15372 8040 -15332 8760
rect -14612 8040 -14572 8760
rect -15372 8000 -14572 8040
rect -13960 8760 -13160 8800
rect -13960 8040 -13920 8760
rect -13200 8040 -13160 8760
rect -13960 8000 -13160 8040
rect -12548 8760 -11748 8800
rect -12548 8040 -12508 8760
rect -11788 8040 -11748 8760
rect -12548 8000 -11748 8040
rect -11136 8760 -10336 8800
rect -11136 8040 -11096 8760
rect -10376 8040 -10336 8760
rect -11136 8000 -10336 8040
rect -9724 8760 -8924 8800
rect -9724 8040 -9684 8760
rect -8964 8040 -8924 8760
rect -9724 8000 -8924 8040
rect -8312 8760 -7512 8800
rect -8312 8040 -8272 8760
rect -7552 8040 -7512 8760
rect -8312 8000 -7512 8040
rect -6900 8760 -6100 8800
rect -6900 8040 -6860 8760
rect -6140 8040 -6100 8760
rect -6900 8000 -6100 8040
rect -5488 8760 -4688 8800
rect -5488 8040 -5448 8760
rect -4728 8040 -4688 8760
rect -5488 8000 -4688 8040
rect -4076 8760 -3276 8800
rect -4076 8040 -4036 8760
rect -3316 8040 -3276 8760
rect -4076 8000 -3276 8040
rect -2664 8760 -1864 8800
rect -2664 8040 -2624 8760
rect -1904 8040 -1864 8760
rect -2664 8000 -1864 8040
rect -1252 8760 -452 8800
rect -1252 8040 -1212 8760
rect -492 8040 -452 8760
rect -1252 8000 -452 8040
rect 160 8760 960 8800
rect 160 8040 200 8760
rect 920 8040 960 8760
rect 160 8000 960 8040
rect 1572 8760 2372 8800
rect 1572 8040 1612 8760
rect 2332 8040 2372 8760
rect 1572 8000 2372 8040
rect 2984 8760 3784 8800
rect 2984 8040 3024 8760
rect 3744 8040 3784 8760
rect 2984 8000 3784 8040
rect 4396 8760 5196 8800
rect 4396 8040 4436 8760
rect 5156 8040 5196 8760
rect 4396 8000 5196 8040
rect 5808 8760 6608 8800
rect 5808 8040 5848 8760
rect 6568 8040 6608 8760
rect 5808 8000 6608 8040
rect 7220 8760 8020 8800
rect 7220 8040 7260 8760
rect 7980 8040 8020 8760
rect 7220 8000 8020 8040
rect 8632 8760 9432 8800
rect 8632 8040 8672 8760
rect 9392 8040 9432 8760
rect 8632 8000 9432 8040
rect 10044 8760 10844 8800
rect 10044 8040 10084 8760
rect 10804 8040 10844 8760
rect 10044 8000 10844 8040
rect 11456 8760 12256 8800
rect 11456 8040 11496 8760
rect 12216 8040 12256 8760
rect 11456 8000 12256 8040
rect 12868 8760 13668 8800
rect 12868 8040 12908 8760
rect 13628 8040 13668 8760
rect 12868 8000 13668 8040
rect 14280 8760 15080 8800
rect 14280 8040 14320 8760
rect 15040 8040 15080 8760
rect 14280 8000 15080 8040
rect 15692 8760 16492 8800
rect 15692 8040 15732 8760
rect 16452 8040 16492 8760
rect 15692 8000 16492 8040
rect 17104 8760 17904 8800
rect 17104 8040 17144 8760
rect 17864 8040 17904 8760
rect 17104 8000 17904 8040
rect 18516 8760 19316 8800
rect 18516 8040 18556 8760
rect 19276 8040 19316 8760
rect 18516 8000 19316 8040
rect 19928 8760 20728 8800
rect 19928 8040 19968 8760
rect 20688 8040 20728 8760
rect 19928 8000 20728 8040
rect 21340 8760 22140 8800
rect 21340 8040 21380 8760
rect 22100 8040 22140 8760
rect 21340 8000 22140 8040
rect 22752 8760 23552 8800
rect 22752 8040 22792 8760
rect 23512 8040 23552 8760
rect 22752 8000 23552 8040
rect -23844 7640 -23044 7680
rect -23844 6920 -23804 7640
rect -23084 6920 -23044 7640
rect -23844 6880 -23044 6920
rect -22432 7640 -21632 7680
rect -22432 6920 -22392 7640
rect -21672 6920 -21632 7640
rect -22432 6880 -21632 6920
rect -21020 7640 -20220 7680
rect -21020 6920 -20980 7640
rect -20260 6920 -20220 7640
rect -21020 6880 -20220 6920
rect -19608 7640 -18808 7680
rect -19608 6920 -19568 7640
rect -18848 6920 -18808 7640
rect -19608 6880 -18808 6920
rect -18196 7640 -17396 7680
rect -18196 6920 -18156 7640
rect -17436 6920 -17396 7640
rect -18196 6880 -17396 6920
rect -16784 7640 -15984 7680
rect -16784 6920 -16744 7640
rect -16024 6920 -15984 7640
rect -16784 6880 -15984 6920
rect -15372 7640 -14572 7680
rect -15372 6920 -15332 7640
rect -14612 6920 -14572 7640
rect -15372 6880 -14572 6920
rect -13960 7640 -13160 7680
rect -13960 6920 -13920 7640
rect -13200 6920 -13160 7640
rect -13960 6880 -13160 6920
rect -12548 7640 -11748 7680
rect -12548 6920 -12508 7640
rect -11788 6920 -11748 7640
rect -12548 6880 -11748 6920
rect -11136 7640 -10336 7680
rect -11136 6920 -11096 7640
rect -10376 6920 -10336 7640
rect -11136 6880 -10336 6920
rect -9724 7640 -8924 7680
rect -9724 6920 -9684 7640
rect -8964 6920 -8924 7640
rect -9724 6880 -8924 6920
rect -8312 7640 -7512 7680
rect -8312 6920 -8272 7640
rect -7552 6920 -7512 7640
rect -8312 6880 -7512 6920
rect -6900 7640 -6100 7680
rect -6900 6920 -6860 7640
rect -6140 6920 -6100 7640
rect -6900 6880 -6100 6920
rect -5488 7640 -4688 7680
rect -5488 6920 -5448 7640
rect -4728 6920 -4688 7640
rect -5488 6880 -4688 6920
rect -4076 7640 -3276 7680
rect -4076 6920 -4036 7640
rect -3316 6920 -3276 7640
rect -4076 6880 -3276 6920
rect -2664 7640 -1864 7680
rect -2664 6920 -2624 7640
rect -1904 6920 -1864 7640
rect -2664 6880 -1864 6920
rect -1252 7640 -452 7680
rect -1252 6920 -1212 7640
rect -492 6920 -452 7640
rect -1252 6880 -452 6920
rect 160 7640 960 7680
rect 160 6920 200 7640
rect 920 6920 960 7640
rect 160 6880 960 6920
rect 1572 7640 2372 7680
rect 1572 6920 1612 7640
rect 2332 6920 2372 7640
rect 1572 6880 2372 6920
rect 2984 7640 3784 7680
rect 2984 6920 3024 7640
rect 3744 6920 3784 7640
rect 2984 6880 3784 6920
rect 4396 7640 5196 7680
rect 4396 6920 4436 7640
rect 5156 6920 5196 7640
rect 4396 6880 5196 6920
rect 5808 7640 6608 7680
rect 5808 6920 5848 7640
rect 6568 6920 6608 7640
rect 5808 6880 6608 6920
rect 7220 7640 8020 7680
rect 7220 6920 7260 7640
rect 7980 6920 8020 7640
rect 7220 6880 8020 6920
rect 8632 7640 9432 7680
rect 8632 6920 8672 7640
rect 9392 6920 9432 7640
rect 8632 6880 9432 6920
rect 10044 7640 10844 7680
rect 10044 6920 10084 7640
rect 10804 6920 10844 7640
rect 10044 6880 10844 6920
rect 11456 7640 12256 7680
rect 11456 6920 11496 7640
rect 12216 6920 12256 7640
rect 11456 6880 12256 6920
rect 12868 7640 13668 7680
rect 12868 6920 12908 7640
rect 13628 6920 13668 7640
rect 12868 6880 13668 6920
rect 14280 7640 15080 7680
rect 14280 6920 14320 7640
rect 15040 6920 15080 7640
rect 14280 6880 15080 6920
rect 15692 7640 16492 7680
rect 15692 6920 15732 7640
rect 16452 6920 16492 7640
rect 15692 6880 16492 6920
rect 17104 7640 17904 7680
rect 17104 6920 17144 7640
rect 17864 6920 17904 7640
rect 17104 6880 17904 6920
rect 18516 7640 19316 7680
rect 18516 6920 18556 7640
rect 19276 6920 19316 7640
rect 18516 6880 19316 6920
rect 19928 7640 20728 7680
rect 19928 6920 19968 7640
rect 20688 6920 20728 7640
rect 19928 6880 20728 6920
rect 21340 7640 22140 7680
rect 21340 6920 21380 7640
rect 22100 6920 22140 7640
rect 21340 6880 22140 6920
rect 22752 7640 23552 7680
rect 22752 6920 22792 7640
rect 23512 6920 23552 7640
rect 22752 6880 23552 6920
rect -23844 6520 -23044 6560
rect -23844 5800 -23804 6520
rect -23084 5800 -23044 6520
rect -23844 5760 -23044 5800
rect -22432 6520 -21632 6560
rect -22432 5800 -22392 6520
rect -21672 5800 -21632 6520
rect -22432 5760 -21632 5800
rect -21020 6520 -20220 6560
rect -21020 5800 -20980 6520
rect -20260 5800 -20220 6520
rect -21020 5760 -20220 5800
rect -19608 6520 -18808 6560
rect -19608 5800 -19568 6520
rect -18848 5800 -18808 6520
rect -19608 5760 -18808 5800
rect -18196 6520 -17396 6560
rect -18196 5800 -18156 6520
rect -17436 5800 -17396 6520
rect -18196 5760 -17396 5800
rect -16784 6520 -15984 6560
rect -16784 5800 -16744 6520
rect -16024 5800 -15984 6520
rect -16784 5760 -15984 5800
rect -15372 6520 -14572 6560
rect -15372 5800 -15332 6520
rect -14612 5800 -14572 6520
rect -15372 5760 -14572 5800
rect -13960 6520 -13160 6560
rect -13960 5800 -13920 6520
rect -13200 5800 -13160 6520
rect -13960 5760 -13160 5800
rect -12548 6520 -11748 6560
rect -12548 5800 -12508 6520
rect -11788 5800 -11748 6520
rect -12548 5760 -11748 5800
rect -11136 6520 -10336 6560
rect -11136 5800 -11096 6520
rect -10376 5800 -10336 6520
rect -11136 5760 -10336 5800
rect -9724 6520 -8924 6560
rect -9724 5800 -9684 6520
rect -8964 5800 -8924 6520
rect -9724 5760 -8924 5800
rect -8312 6520 -7512 6560
rect -8312 5800 -8272 6520
rect -7552 5800 -7512 6520
rect -8312 5760 -7512 5800
rect -6900 6520 -6100 6560
rect -6900 5800 -6860 6520
rect -6140 5800 -6100 6520
rect -6900 5760 -6100 5800
rect -5488 6520 -4688 6560
rect -5488 5800 -5448 6520
rect -4728 5800 -4688 6520
rect -5488 5760 -4688 5800
rect -4076 6520 -3276 6560
rect -4076 5800 -4036 6520
rect -3316 5800 -3276 6520
rect -4076 5760 -3276 5800
rect -2664 6520 -1864 6560
rect -2664 5800 -2624 6520
rect -1904 5800 -1864 6520
rect -2664 5760 -1864 5800
rect -1252 6520 -452 6560
rect -1252 5800 -1212 6520
rect -492 5800 -452 6520
rect -1252 5760 -452 5800
rect 160 6520 960 6560
rect 160 5800 200 6520
rect 920 5800 960 6520
rect 160 5760 960 5800
rect 1572 6520 2372 6560
rect 1572 5800 1612 6520
rect 2332 5800 2372 6520
rect 1572 5760 2372 5800
rect 2984 6520 3784 6560
rect 2984 5800 3024 6520
rect 3744 5800 3784 6520
rect 2984 5760 3784 5800
rect 4396 6520 5196 6560
rect 4396 5800 4436 6520
rect 5156 5800 5196 6520
rect 4396 5760 5196 5800
rect 5808 6520 6608 6560
rect 5808 5800 5848 6520
rect 6568 5800 6608 6520
rect 5808 5760 6608 5800
rect 7220 6520 8020 6560
rect 7220 5800 7260 6520
rect 7980 5800 8020 6520
rect 7220 5760 8020 5800
rect 8632 6520 9432 6560
rect 8632 5800 8672 6520
rect 9392 5800 9432 6520
rect 8632 5760 9432 5800
rect 10044 6520 10844 6560
rect 10044 5800 10084 6520
rect 10804 5800 10844 6520
rect 10044 5760 10844 5800
rect 11456 6520 12256 6560
rect 11456 5800 11496 6520
rect 12216 5800 12256 6520
rect 11456 5760 12256 5800
rect 12868 6520 13668 6560
rect 12868 5800 12908 6520
rect 13628 5800 13668 6520
rect 12868 5760 13668 5800
rect 14280 6520 15080 6560
rect 14280 5800 14320 6520
rect 15040 5800 15080 6520
rect 14280 5760 15080 5800
rect 15692 6520 16492 6560
rect 15692 5800 15732 6520
rect 16452 5800 16492 6520
rect 15692 5760 16492 5800
rect 17104 6520 17904 6560
rect 17104 5800 17144 6520
rect 17864 5800 17904 6520
rect 17104 5760 17904 5800
rect 18516 6520 19316 6560
rect 18516 5800 18556 6520
rect 19276 5800 19316 6520
rect 18516 5760 19316 5800
rect 19928 6520 20728 6560
rect 19928 5800 19968 6520
rect 20688 5800 20728 6520
rect 19928 5760 20728 5800
rect 21340 6520 22140 6560
rect 21340 5800 21380 6520
rect 22100 5800 22140 6520
rect 21340 5760 22140 5800
rect 22752 6520 23552 6560
rect 22752 5800 22792 6520
rect 23512 5800 23552 6520
rect 22752 5760 23552 5800
rect -23844 5400 -23044 5440
rect -23844 4680 -23804 5400
rect -23084 4680 -23044 5400
rect -23844 4640 -23044 4680
rect -22432 5400 -21632 5440
rect -22432 4680 -22392 5400
rect -21672 4680 -21632 5400
rect -22432 4640 -21632 4680
rect -21020 5400 -20220 5440
rect -21020 4680 -20980 5400
rect -20260 4680 -20220 5400
rect -21020 4640 -20220 4680
rect -19608 5400 -18808 5440
rect -19608 4680 -19568 5400
rect -18848 4680 -18808 5400
rect -19608 4640 -18808 4680
rect -18196 5400 -17396 5440
rect -18196 4680 -18156 5400
rect -17436 4680 -17396 5400
rect -18196 4640 -17396 4680
rect -16784 5400 -15984 5440
rect -16784 4680 -16744 5400
rect -16024 4680 -15984 5400
rect -16784 4640 -15984 4680
rect -15372 5400 -14572 5440
rect -15372 4680 -15332 5400
rect -14612 4680 -14572 5400
rect -15372 4640 -14572 4680
rect -13960 5400 -13160 5440
rect -13960 4680 -13920 5400
rect -13200 4680 -13160 5400
rect -13960 4640 -13160 4680
rect -12548 5400 -11748 5440
rect -12548 4680 -12508 5400
rect -11788 4680 -11748 5400
rect -12548 4640 -11748 4680
rect -11136 5400 -10336 5440
rect -11136 4680 -11096 5400
rect -10376 4680 -10336 5400
rect -11136 4640 -10336 4680
rect -9724 5400 -8924 5440
rect -9724 4680 -9684 5400
rect -8964 4680 -8924 5400
rect -9724 4640 -8924 4680
rect -8312 5400 -7512 5440
rect -8312 4680 -8272 5400
rect -7552 4680 -7512 5400
rect -8312 4640 -7512 4680
rect -6900 5400 -6100 5440
rect -6900 4680 -6860 5400
rect -6140 4680 -6100 5400
rect -6900 4640 -6100 4680
rect -5488 5400 -4688 5440
rect -5488 4680 -5448 5400
rect -4728 4680 -4688 5400
rect -5488 4640 -4688 4680
rect -4076 5400 -3276 5440
rect -4076 4680 -4036 5400
rect -3316 4680 -3276 5400
rect -4076 4640 -3276 4680
rect -2664 5400 -1864 5440
rect -2664 4680 -2624 5400
rect -1904 4680 -1864 5400
rect -2664 4640 -1864 4680
rect -1252 5400 -452 5440
rect -1252 4680 -1212 5400
rect -492 4680 -452 5400
rect -1252 4640 -452 4680
rect 160 5400 960 5440
rect 160 4680 200 5400
rect 920 4680 960 5400
rect 160 4640 960 4680
rect 1572 5400 2372 5440
rect 1572 4680 1612 5400
rect 2332 4680 2372 5400
rect 1572 4640 2372 4680
rect 2984 5400 3784 5440
rect 2984 4680 3024 5400
rect 3744 4680 3784 5400
rect 2984 4640 3784 4680
rect 4396 5400 5196 5440
rect 4396 4680 4436 5400
rect 5156 4680 5196 5400
rect 4396 4640 5196 4680
rect 5808 5400 6608 5440
rect 5808 4680 5848 5400
rect 6568 4680 6608 5400
rect 5808 4640 6608 4680
rect 7220 5400 8020 5440
rect 7220 4680 7260 5400
rect 7980 4680 8020 5400
rect 7220 4640 8020 4680
rect 8632 5400 9432 5440
rect 8632 4680 8672 5400
rect 9392 4680 9432 5400
rect 8632 4640 9432 4680
rect 10044 5400 10844 5440
rect 10044 4680 10084 5400
rect 10804 4680 10844 5400
rect 10044 4640 10844 4680
rect 11456 5400 12256 5440
rect 11456 4680 11496 5400
rect 12216 4680 12256 5400
rect 11456 4640 12256 4680
rect 12868 5400 13668 5440
rect 12868 4680 12908 5400
rect 13628 4680 13668 5400
rect 12868 4640 13668 4680
rect 14280 5400 15080 5440
rect 14280 4680 14320 5400
rect 15040 4680 15080 5400
rect 14280 4640 15080 4680
rect 15692 5400 16492 5440
rect 15692 4680 15732 5400
rect 16452 4680 16492 5400
rect 15692 4640 16492 4680
rect 17104 5400 17904 5440
rect 17104 4680 17144 5400
rect 17864 4680 17904 5400
rect 17104 4640 17904 4680
rect 18516 5400 19316 5440
rect 18516 4680 18556 5400
rect 19276 4680 19316 5400
rect 18516 4640 19316 4680
rect 19928 5400 20728 5440
rect 19928 4680 19968 5400
rect 20688 4680 20728 5400
rect 19928 4640 20728 4680
rect 21340 5400 22140 5440
rect 21340 4680 21380 5400
rect 22100 4680 22140 5400
rect 21340 4640 22140 4680
rect 22752 5400 23552 5440
rect 22752 4680 22792 5400
rect 23512 4680 23552 5400
rect 22752 4640 23552 4680
rect -23844 4280 -23044 4320
rect -23844 3560 -23804 4280
rect -23084 3560 -23044 4280
rect -23844 3520 -23044 3560
rect -22432 4280 -21632 4320
rect -22432 3560 -22392 4280
rect -21672 3560 -21632 4280
rect -22432 3520 -21632 3560
rect -21020 4280 -20220 4320
rect -21020 3560 -20980 4280
rect -20260 3560 -20220 4280
rect -21020 3520 -20220 3560
rect -19608 4280 -18808 4320
rect -19608 3560 -19568 4280
rect -18848 3560 -18808 4280
rect -19608 3520 -18808 3560
rect -18196 4280 -17396 4320
rect -18196 3560 -18156 4280
rect -17436 3560 -17396 4280
rect -18196 3520 -17396 3560
rect -16784 4280 -15984 4320
rect -16784 3560 -16744 4280
rect -16024 3560 -15984 4280
rect -16784 3520 -15984 3560
rect -15372 4280 -14572 4320
rect -15372 3560 -15332 4280
rect -14612 3560 -14572 4280
rect -15372 3520 -14572 3560
rect -13960 4280 -13160 4320
rect -13960 3560 -13920 4280
rect -13200 3560 -13160 4280
rect -13960 3520 -13160 3560
rect -12548 4280 -11748 4320
rect -12548 3560 -12508 4280
rect -11788 3560 -11748 4280
rect -12548 3520 -11748 3560
rect -11136 4280 -10336 4320
rect -11136 3560 -11096 4280
rect -10376 3560 -10336 4280
rect -11136 3520 -10336 3560
rect -9724 4280 -8924 4320
rect -9724 3560 -9684 4280
rect -8964 3560 -8924 4280
rect -9724 3520 -8924 3560
rect -8312 4280 -7512 4320
rect -8312 3560 -8272 4280
rect -7552 3560 -7512 4280
rect -8312 3520 -7512 3560
rect -6900 4280 -6100 4320
rect -6900 3560 -6860 4280
rect -6140 3560 -6100 4280
rect -6900 3520 -6100 3560
rect -5488 4280 -4688 4320
rect -5488 3560 -5448 4280
rect -4728 3560 -4688 4280
rect -5488 3520 -4688 3560
rect -4076 4280 -3276 4320
rect -4076 3560 -4036 4280
rect -3316 3560 -3276 4280
rect -4076 3520 -3276 3560
rect -2664 4280 -1864 4320
rect -2664 3560 -2624 4280
rect -1904 3560 -1864 4280
rect -2664 3520 -1864 3560
rect -1252 4280 -452 4320
rect -1252 3560 -1212 4280
rect -492 3560 -452 4280
rect -1252 3520 -452 3560
rect 160 4280 960 4320
rect 160 3560 200 4280
rect 920 3560 960 4280
rect 160 3520 960 3560
rect 1572 4280 2372 4320
rect 1572 3560 1612 4280
rect 2332 3560 2372 4280
rect 1572 3520 2372 3560
rect 2984 4280 3784 4320
rect 2984 3560 3024 4280
rect 3744 3560 3784 4280
rect 2984 3520 3784 3560
rect 4396 4280 5196 4320
rect 4396 3560 4436 4280
rect 5156 3560 5196 4280
rect 4396 3520 5196 3560
rect 5808 4280 6608 4320
rect 5808 3560 5848 4280
rect 6568 3560 6608 4280
rect 5808 3520 6608 3560
rect 7220 4280 8020 4320
rect 7220 3560 7260 4280
rect 7980 3560 8020 4280
rect 7220 3520 8020 3560
rect 8632 4280 9432 4320
rect 8632 3560 8672 4280
rect 9392 3560 9432 4280
rect 8632 3520 9432 3560
rect 10044 4280 10844 4320
rect 10044 3560 10084 4280
rect 10804 3560 10844 4280
rect 10044 3520 10844 3560
rect 11456 4280 12256 4320
rect 11456 3560 11496 4280
rect 12216 3560 12256 4280
rect 11456 3520 12256 3560
rect 12868 4280 13668 4320
rect 12868 3560 12908 4280
rect 13628 3560 13668 4280
rect 12868 3520 13668 3560
rect 14280 4280 15080 4320
rect 14280 3560 14320 4280
rect 15040 3560 15080 4280
rect 14280 3520 15080 3560
rect 15692 4280 16492 4320
rect 15692 3560 15732 4280
rect 16452 3560 16492 4280
rect 15692 3520 16492 3560
rect 17104 4280 17904 4320
rect 17104 3560 17144 4280
rect 17864 3560 17904 4280
rect 17104 3520 17904 3560
rect 18516 4280 19316 4320
rect 18516 3560 18556 4280
rect 19276 3560 19316 4280
rect 18516 3520 19316 3560
rect 19928 4280 20728 4320
rect 19928 3560 19968 4280
rect 20688 3560 20728 4280
rect 19928 3520 20728 3560
rect 21340 4280 22140 4320
rect 21340 3560 21380 4280
rect 22100 3560 22140 4280
rect 21340 3520 22140 3560
rect 22752 4280 23552 4320
rect 22752 3560 22792 4280
rect 23512 3560 23552 4280
rect 22752 3520 23552 3560
rect -23844 3160 -23044 3200
rect -23844 2440 -23804 3160
rect -23084 2440 -23044 3160
rect -23844 2400 -23044 2440
rect -22432 3160 -21632 3200
rect -22432 2440 -22392 3160
rect -21672 2440 -21632 3160
rect -22432 2400 -21632 2440
rect -21020 3160 -20220 3200
rect -21020 2440 -20980 3160
rect -20260 2440 -20220 3160
rect -21020 2400 -20220 2440
rect -19608 3160 -18808 3200
rect -19608 2440 -19568 3160
rect -18848 2440 -18808 3160
rect -19608 2400 -18808 2440
rect -18196 3160 -17396 3200
rect -18196 2440 -18156 3160
rect -17436 2440 -17396 3160
rect -18196 2400 -17396 2440
rect -16784 3160 -15984 3200
rect -16784 2440 -16744 3160
rect -16024 2440 -15984 3160
rect -16784 2400 -15984 2440
rect -15372 3160 -14572 3200
rect -15372 2440 -15332 3160
rect -14612 2440 -14572 3160
rect -15372 2400 -14572 2440
rect -13960 3160 -13160 3200
rect -13960 2440 -13920 3160
rect -13200 2440 -13160 3160
rect -13960 2400 -13160 2440
rect -12548 3160 -11748 3200
rect -12548 2440 -12508 3160
rect -11788 2440 -11748 3160
rect -12548 2400 -11748 2440
rect -11136 3160 -10336 3200
rect -11136 2440 -11096 3160
rect -10376 2440 -10336 3160
rect -11136 2400 -10336 2440
rect -9724 3160 -8924 3200
rect -9724 2440 -9684 3160
rect -8964 2440 -8924 3160
rect -9724 2400 -8924 2440
rect -8312 3160 -7512 3200
rect -8312 2440 -8272 3160
rect -7552 2440 -7512 3160
rect -8312 2400 -7512 2440
rect -6900 3160 -6100 3200
rect -6900 2440 -6860 3160
rect -6140 2440 -6100 3160
rect -6900 2400 -6100 2440
rect -5488 3160 -4688 3200
rect -5488 2440 -5448 3160
rect -4728 2440 -4688 3160
rect -5488 2400 -4688 2440
rect -4076 3160 -3276 3200
rect -4076 2440 -4036 3160
rect -3316 2440 -3276 3160
rect -4076 2400 -3276 2440
rect -2664 3160 -1864 3200
rect -2664 2440 -2624 3160
rect -1904 2440 -1864 3160
rect -2664 2400 -1864 2440
rect -1252 3160 -452 3200
rect -1252 2440 -1212 3160
rect -492 2440 -452 3160
rect -1252 2400 -452 2440
rect 160 3160 960 3200
rect 160 2440 200 3160
rect 920 2440 960 3160
rect 160 2400 960 2440
rect 1572 3160 2372 3200
rect 1572 2440 1612 3160
rect 2332 2440 2372 3160
rect 1572 2400 2372 2440
rect 2984 3160 3784 3200
rect 2984 2440 3024 3160
rect 3744 2440 3784 3160
rect 2984 2400 3784 2440
rect 4396 3160 5196 3200
rect 4396 2440 4436 3160
rect 5156 2440 5196 3160
rect 4396 2400 5196 2440
rect 5808 3160 6608 3200
rect 5808 2440 5848 3160
rect 6568 2440 6608 3160
rect 5808 2400 6608 2440
rect 7220 3160 8020 3200
rect 7220 2440 7260 3160
rect 7980 2440 8020 3160
rect 7220 2400 8020 2440
rect 8632 3160 9432 3200
rect 8632 2440 8672 3160
rect 9392 2440 9432 3160
rect 8632 2400 9432 2440
rect 10044 3160 10844 3200
rect 10044 2440 10084 3160
rect 10804 2440 10844 3160
rect 10044 2400 10844 2440
rect 11456 3160 12256 3200
rect 11456 2440 11496 3160
rect 12216 2440 12256 3160
rect 11456 2400 12256 2440
rect 12868 3160 13668 3200
rect 12868 2440 12908 3160
rect 13628 2440 13668 3160
rect 12868 2400 13668 2440
rect 14280 3160 15080 3200
rect 14280 2440 14320 3160
rect 15040 2440 15080 3160
rect 14280 2400 15080 2440
rect 15692 3160 16492 3200
rect 15692 2440 15732 3160
rect 16452 2440 16492 3160
rect 15692 2400 16492 2440
rect 17104 3160 17904 3200
rect 17104 2440 17144 3160
rect 17864 2440 17904 3160
rect 17104 2400 17904 2440
rect 18516 3160 19316 3200
rect 18516 2440 18556 3160
rect 19276 2440 19316 3160
rect 18516 2400 19316 2440
rect 19928 3160 20728 3200
rect 19928 2440 19968 3160
rect 20688 2440 20728 3160
rect 19928 2400 20728 2440
rect 21340 3160 22140 3200
rect 21340 2440 21380 3160
rect 22100 2440 22140 3160
rect 21340 2400 22140 2440
rect 22752 3160 23552 3200
rect 22752 2440 22792 3160
rect 23512 2440 23552 3160
rect 22752 2400 23552 2440
rect -23844 2040 -23044 2080
rect -23844 1320 -23804 2040
rect -23084 1320 -23044 2040
rect -23844 1280 -23044 1320
rect -22432 2040 -21632 2080
rect -22432 1320 -22392 2040
rect -21672 1320 -21632 2040
rect -22432 1280 -21632 1320
rect -21020 2040 -20220 2080
rect -21020 1320 -20980 2040
rect -20260 1320 -20220 2040
rect -21020 1280 -20220 1320
rect -19608 2040 -18808 2080
rect -19608 1320 -19568 2040
rect -18848 1320 -18808 2040
rect -19608 1280 -18808 1320
rect -18196 2040 -17396 2080
rect -18196 1320 -18156 2040
rect -17436 1320 -17396 2040
rect -18196 1280 -17396 1320
rect -16784 2040 -15984 2080
rect -16784 1320 -16744 2040
rect -16024 1320 -15984 2040
rect -16784 1280 -15984 1320
rect -15372 2040 -14572 2080
rect -15372 1320 -15332 2040
rect -14612 1320 -14572 2040
rect -15372 1280 -14572 1320
rect -13960 2040 -13160 2080
rect -13960 1320 -13920 2040
rect -13200 1320 -13160 2040
rect -13960 1280 -13160 1320
rect -12548 2040 -11748 2080
rect -12548 1320 -12508 2040
rect -11788 1320 -11748 2040
rect -12548 1280 -11748 1320
rect -11136 2040 -10336 2080
rect -11136 1320 -11096 2040
rect -10376 1320 -10336 2040
rect -11136 1280 -10336 1320
rect -9724 2040 -8924 2080
rect -9724 1320 -9684 2040
rect -8964 1320 -8924 2040
rect -9724 1280 -8924 1320
rect -8312 2040 -7512 2080
rect -8312 1320 -8272 2040
rect -7552 1320 -7512 2040
rect -8312 1280 -7512 1320
rect -6900 2040 -6100 2080
rect -6900 1320 -6860 2040
rect -6140 1320 -6100 2040
rect -6900 1280 -6100 1320
rect -5488 2040 -4688 2080
rect -5488 1320 -5448 2040
rect -4728 1320 -4688 2040
rect -5488 1280 -4688 1320
rect -4076 2040 -3276 2080
rect -4076 1320 -4036 2040
rect -3316 1320 -3276 2040
rect -4076 1280 -3276 1320
rect -2664 2040 -1864 2080
rect -2664 1320 -2624 2040
rect -1904 1320 -1864 2040
rect -2664 1280 -1864 1320
rect -1252 2040 -452 2080
rect -1252 1320 -1212 2040
rect -492 1320 -452 2040
rect -1252 1280 -452 1320
rect 160 2040 960 2080
rect 160 1320 200 2040
rect 920 1320 960 2040
rect 160 1280 960 1320
rect 1572 2040 2372 2080
rect 1572 1320 1612 2040
rect 2332 1320 2372 2040
rect 1572 1280 2372 1320
rect 2984 2040 3784 2080
rect 2984 1320 3024 2040
rect 3744 1320 3784 2040
rect 2984 1280 3784 1320
rect 4396 2040 5196 2080
rect 4396 1320 4436 2040
rect 5156 1320 5196 2040
rect 4396 1280 5196 1320
rect 5808 2040 6608 2080
rect 5808 1320 5848 2040
rect 6568 1320 6608 2040
rect 5808 1280 6608 1320
rect 7220 2040 8020 2080
rect 7220 1320 7260 2040
rect 7980 1320 8020 2040
rect 7220 1280 8020 1320
rect 8632 2040 9432 2080
rect 8632 1320 8672 2040
rect 9392 1320 9432 2040
rect 8632 1280 9432 1320
rect 10044 2040 10844 2080
rect 10044 1320 10084 2040
rect 10804 1320 10844 2040
rect 10044 1280 10844 1320
rect 11456 2040 12256 2080
rect 11456 1320 11496 2040
rect 12216 1320 12256 2040
rect 11456 1280 12256 1320
rect 12868 2040 13668 2080
rect 12868 1320 12908 2040
rect 13628 1320 13668 2040
rect 12868 1280 13668 1320
rect 14280 2040 15080 2080
rect 14280 1320 14320 2040
rect 15040 1320 15080 2040
rect 14280 1280 15080 1320
rect 15692 2040 16492 2080
rect 15692 1320 15732 2040
rect 16452 1320 16492 2040
rect 15692 1280 16492 1320
rect 17104 2040 17904 2080
rect 17104 1320 17144 2040
rect 17864 1320 17904 2040
rect 17104 1280 17904 1320
rect 18516 2040 19316 2080
rect 18516 1320 18556 2040
rect 19276 1320 19316 2040
rect 18516 1280 19316 1320
rect 19928 2040 20728 2080
rect 19928 1320 19968 2040
rect 20688 1320 20728 2040
rect 19928 1280 20728 1320
rect 21340 2040 22140 2080
rect 21340 1320 21380 2040
rect 22100 1320 22140 2040
rect 21340 1280 22140 1320
rect 22752 2040 23552 2080
rect 22752 1320 22792 2040
rect 23512 1320 23552 2040
rect 22752 1280 23552 1320
rect -23844 920 -23044 960
rect -23844 200 -23804 920
rect -23084 200 -23044 920
rect -23844 160 -23044 200
rect -22432 920 -21632 960
rect -22432 200 -22392 920
rect -21672 200 -21632 920
rect -22432 160 -21632 200
rect -21020 920 -20220 960
rect -21020 200 -20980 920
rect -20260 200 -20220 920
rect -21020 160 -20220 200
rect -19608 920 -18808 960
rect -19608 200 -19568 920
rect -18848 200 -18808 920
rect -19608 160 -18808 200
rect -18196 920 -17396 960
rect -18196 200 -18156 920
rect -17436 200 -17396 920
rect -18196 160 -17396 200
rect -16784 920 -15984 960
rect -16784 200 -16744 920
rect -16024 200 -15984 920
rect -16784 160 -15984 200
rect -15372 920 -14572 960
rect -15372 200 -15332 920
rect -14612 200 -14572 920
rect -15372 160 -14572 200
rect -13960 920 -13160 960
rect -13960 200 -13920 920
rect -13200 200 -13160 920
rect -13960 160 -13160 200
rect -12548 920 -11748 960
rect -12548 200 -12508 920
rect -11788 200 -11748 920
rect -12548 160 -11748 200
rect -11136 920 -10336 960
rect -11136 200 -11096 920
rect -10376 200 -10336 920
rect -11136 160 -10336 200
rect -9724 920 -8924 960
rect -9724 200 -9684 920
rect -8964 200 -8924 920
rect -9724 160 -8924 200
rect -8312 920 -7512 960
rect -8312 200 -8272 920
rect -7552 200 -7512 920
rect -8312 160 -7512 200
rect -6900 920 -6100 960
rect -6900 200 -6860 920
rect -6140 200 -6100 920
rect -6900 160 -6100 200
rect -5488 920 -4688 960
rect -5488 200 -5448 920
rect -4728 200 -4688 920
rect -5488 160 -4688 200
rect -4076 920 -3276 960
rect -4076 200 -4036 920
rect -3316 200 -3276 920
rect -4076 160 -3276 200
rect -2664 920 -1864 960
rect -2664 200 -2624 920
rect -1904 200 -1864 920
rect -2664 160 -1864 200
rect -1252 920 -452 960
rect -1252 200 -1212 920
rect -492 200 -452 920
rect -1252 160 -452 200
rect 160 920 960 960
rect 160 200 200 920
rect 920 200 960 920
rect 160 160 960 200
rect 1572 920 2372 960
rect 1572 200 1612 920
rect 2332 200 2372 920
rect 1572 160 2372 200
rect 2984 920 3784 960
rect 2984 200 3024 920
rect 3744 200 3784 920
rect 2984 160 3784 200
rect 4396 920 5196 960
rect 4396 200 4436 920
rect 5156 200 5196 920
rect 4396 160 5196 200
rect 5808 920 6608 960
rect 5808 200 5848 920
rect 6568 200 6608 920
rect 5808 160 6608 200
rect 7220 920 8020 960
rect 7220 200 7260 920
rect 7980 200 8020 920
rect 7220 160 8020 200
rect 8632 920 9432 960
rect 8632 200 8672 920
rect 9392 200 9432 920
rect 8632 160 9432 200
rect 10044 920 10844 960
rect 10044 200 10084 920
rect 10804 200 10844 920
rect 10044 160 10844 200
rect 11456 920 12256 960
rect 11456 200 11496 920
rect 12216 200 12256 920
rect 11456 160 12256 200
rect 12868 920 13668 960
rect 12868 200 12908 920
rect 13628 200 13668 920
rect 12868 160 13668 200
rect 14280 920 15080 960
rect 14280 200 14320 920
rect 15040 200 15080 920
rect 14280 160 15080 200
rect 15692 920 16492 960
rect 15692 200 15732 920
rect 16452 200 16492 920
rect 15692 160 16492 200
rect 17104 920 17904 960
rect 17104 200 17144 920
rect 17864 200 17904 920
rect 17104 160 17904 200
rect 18516 920 19316 960
rect 18516 200 18556 920
rect 19276 200 19316 920
rect 18516 160 19316 200
rect 19928 920 20728 960
rect 19928 200 19968 920
rect 20688 200 20728 920
rect 19928 160 20728 200
rect 21340 920 22140 960
rect 21340 200 21380 920
rect 22100 200 22140 920
rect 21340 160 22140 200
rect 22752 920 23552 960
rect 22752 200 22792 920
rect 23512 200 23552 920
rect 22752 160 23552 200
rect -23844 -200 -23044 -160
rect -23844 -920 -23804 -200
rect -23084 -920 -23044 -200
rect -23844 -960 -23044 -920
rect -22432 -200 -21632 -160
rect -22432 -920 -22392 -200
rect -21672 -920 -21632 -200
rect -22432 -960 -21632 -920
rect -21020 -200 -20220 -160
rect -21020 -920 -20980 -200
rect -20260 -920 -20220 -200
rect -21020 -960 -20220 -920
rect -19608 -200 -18808 -160
rect -19608 -920 -19568 -200
rect -18848 -920 -18808 -200
rect -19608 -960 -18808 -920
rect -18196 -200 -17396 -160
rect -18196 -920 -18156 -200
rect -17436 -920 -17396 -200
rect -18196 -960 -17396 -920
rect -16784 -200 -15984 -160
rect -16784 -920 -16744 -200
rect -16024 -920 -15984 -200
rect -16784 -960 -15984 -920
rect -15372 -200 -14572 -160
rect -15372 -920 -15332 -200
rect -14612 -920 -14572 -200
rect -15372 -960 -14572 -920
rect -13960 -200 -13160 -160
rect -13960 -920 -13920 -200
rect -13200 -920 -13160 -200
rect -13960 -960 -13160 -920
rect -12548 -200 -11748 -160
rect -12548 -920 -12508 -200
rect -11788 -920 -11748 -200
rect -12548 -960 -11748 -920
rect -11136 -200 -10336 -160
rect -11136 -920 -11096 -200
rect -10376 -920 -10336 -200
rect -11136 -960 -10336 -920
rect -9724 -200 -8924 -160
rect -9724 -920 -9684 -200
rect -8964 -920 -8924 -200
rect -9724 -960 -8924 -920
rect -8312 -200 -7512 -160
rect -8312 -920 -8272 -200
rect -7552 -920 -7512 -200
rect -8312 -960 -7512 -920
rect -6900 -200 -6100 -160
rect -6900 -920 -6860 -200
rect -6140 -920 -6100 -200
rect -6900 -960 -6100 -920
rect -5488 -200 -4688 -160
rect -5488 -920 -5448 -200
rect -4728 -920 -4688 -200
rect -5488 -960 -4688 -920
rect -4076 -200 -3276 -160
rect -4076 -920 -4036 -200
rect -3316 -920 -3276 -200
rect -4076 -960 -3276 -920
rect -2664 -200 -1864 -160
rect -2664 -920 -2624 -200
rect -1904 -920 -1864 -200
rect -2664 -960 -1864 -920
rect -1252 -200 -452 -160
rect -1252 -920 -1212 -200
rect -492 -920 -452 -200
rect -1252 -960 -452 -920
rect 160 -200 960 -160
rect 160 -920 200 -200
rect 920 -920 960 -200
rect 160 -960 960 -920
rect 1572 -200 2372 -160
rect 1572 -920 1612 -200
rect 2332 -920 2372 -200
rect 1572 -960 2372 -920
rect 2984 -200 3784 -160
rect 2984 -920 3024 -200
rect 3744 -920 3784 -200
rect 2984 -960 3784 -920
rect 4396 -200 5196 -160
rect 4396 -920 4436 -200
rect 5156 -920 5196 -200
rect 4396 -960 5196 -920
rect 5808 -200 6608 -160
rect 5808 -920 5848 -200
rect 6568 -920 6608 -200
rect 5808 -960 6608 -920
rect 7220 -200 8020 -160
rect 7220 -920 7260 -200
rect 7980 -920 8020 -200
rect 7220 -960 8020 -920
rect 8632 -200 9432 -160
rect 8632 -920 8672 -200
rect 9392 -920 9432 -200
rect 8632 -960 9432 -920
rect 10044 -200 10844 -160
rect 10044 -920 10084 -200
rect 10804 -920 10844 -200
rect 10044 -960 10844 -920
rect 11456 -200 12256 -160
rect 11456 -920 11496 -200
rect 12216 -920 12256 -200
rect 11456 -960 12256 -920
rect 12868 -200 13668 -160
rect 12868 -920 12908 -200
rect 13628 -920 13668 -200
rect 12868 -960 13668 -920
rect 14280 -200 15080 -160
rect 14280 -920 14320 -200
rect 15040 -920 15080 -200
rect 14280 -960 15080 -920
rect 15692 -200 16492 -160
rect 15692 -920 15732 -200
rect 16452 -920 16492 -200
rect 15692 -960 16492 -920
rect 17104 -200 17904 -160
rect 17104 -920 17144 -200
rect 17864 -920 17904 -200
rect 17104 -960 17904 -920
rect 18516 -200 19316 -160
rect 18516 -920 18556 -200
rect 19276 -920 19316 -200
rect 18516 -960 19316 -920
rect 19928 -200 20728 -160
rect 19928 -920 19968 -200
rect 20688 -920 20728 -200
rect 19928 -960 20728 -920
rect 21340 -200 22140 -160
rect 21340 -920 21380 -200
rect 22100 -920 22140 -200
rect 21340 -960 22140 -920
rect 22752 -200 23552 -160
rect 22752 -920 22792 -200
rect 23512 -920 23552 -200
rect 22752 -960 23552 -920
rect -23844 -1320 -23044 -1280
rect -23844 -2040 -23804 -1320
rect -23084 -2040 -23044 -1320
rect -23844 -2080 -23044 -2040
rect -22432 -1320 -21632 -1280
rect -22432 -2040 -22392 -1320
rect -21672 -2040 -21632 -1320
rect -22432 -2080 -21632 -2040
rect -21020 -1320 -20220 -1280
rect -21020 -2040 -20980 -1320
rect -20260 -2040 -20220 -1320
rect -21020 -2080 -20220 -2040
rect -19608 -1320 -18808 -1280
rect -19608 -2040 -19568 -1320
rect -18848 -2040 -18808 -1320
rect -19608 -2080 -18808 -2040
rect -18196 -1320 -17396 -1280
rect -18196 -2040 -18156 -1320
rect -17436 -2040 -17396 -1320
rect -18196 -2080 -17396 -2040
rect -16784 -1320 -15984 -1280
rect -16784 -2040 -16744 -1320
rect -16024 -2040 -15984 -1320
rect -16784 -2080 -15984 -2040
rect -15372 -1320 -14572 -1280
rect -15372 -2040 -15332 -1320
rect -14612 -2040 -14572 -1320
rect -15372 -2080 -14572 -2040
rect -13960 -1320 -13160 -1280
rect -13960 -2040 -13920 -1320
rect -13200 -2040 -13160 -1320
rect -13960 -2080 -13160 -2040
rect -12548 -1320 -11748 -1280
rect -12548 -2040 -12508 -1320
rect -11788 -2040 -11748 -1320
rect -12548 -2080 -11748 -2040
rect -11136 -1320 -10336 -1280
rect -11136 -2040 -11096 -1320
rect -10376 -2040 -10336 -1320
rect -11136 -2080 -10336 -2040
rect -9724 -1320 -8924 -1280
rect -9724 -2040 -9684 -1320
rect -8964 -2040 -8924 -1320
rect -9724 -2080 -8924 -2040
rect -8312 -1320 -7512 -1280
rect -8312 -2040 -8272 -1320
rect -7552 -2040 -7512 -1320
rect -8312 -2080 -7512 -2040
rect -6900 -1320 -6100 -1280
rect -6900 -2040 -6860 -1320
rect -6140 -2040 -6100 -1320
rect -6900 -2080 -6100 -2040
rect -5488 -1320 -4688 -1280
rect -5488 -2040 -5448 -1320
rect -4728 -2040 -4688 -1320
rect -5488 -2080 -4688 -2040
rect -4076 -1320 -3276 -1280
rect -4076 -2040 -4036 -1320
rect -3316 -2040 -3276 -1320
rect -4076 -2080 -3276 -2040
rect -2664 -1320 -1864 -1280
rect -2664 -2040 -2624 -1320
rect -1904 -2040 -1864 -1320
rect -2664 -2080 -1864 -2040
rect -1252 -1320 -452 -1280
rect -1252 -2040 -1212 -1320
rect -492 -2040 -452 -1320
rect -1252 -2080 -452 -2040
rect 160 -1320 960 -1280
rect 160 -2040 200 -1320
rect 920 -2040 960 -1320
rect 160 -2080 960 -2040
rect 1572 -1320 2372 -1280
rect 1572 -2040 1612 -1320
rect 2332 -2040 2372 -1320
rect 1572 -2080 2372 -2040
rect 2984 -1320 3784 -1280
rect 2984 -2040 3024 -1320
rect 3744 -2040 3784 -1320
rect 2984 -2080 3784 -2040
rect 4396 -1320 5196 -1280
rect 4396 -2040 4436 -1320
rect 5156 -2040 5196 -1320
rect 4396 -2080 5196 -2040
rect 5808 -1320 6608 -1280
rect 5808 -2040 5848 -1320
rect 6568 -2040 6608 -1320
rect 5808 -2080 6608 -2040
rect 7220 -1320 8020 -1280
rect 7220 -2040 7260 -1320
rect 7980 -2040 8020 -1320
rect 7220 -2080 8020 -2040
rect 8632 -1320 9432 -1280
rect 8632 -2040 8672 -1320
rect 9392 -2040 9432 -1320
rect 8632 -2080 9432 -2040
rect 10044 -1320 10844 -1280
rect 10044 -2040 10084 -1320
rect 10804 -2040 10844 -1320
rect 10044 -2080 10844 -2040
rect 11456 -1320 12256 -1280
rect 11456 -2040 11496 -1320
rect 12216 -2040 12256 -1320
rect 11456 -2080 12256 -2040
rect 12868 -1320 13668 -1280
rect 12868 -2040 12908 -1320
rect 13628 -2040 13668 -1320
rect 12868 -2080 13668 -2040
rect 14280 -1320 15080 -1280
rect 14280 -2040 14320 -1320
rect 15040 -2040 15080 -1320
rect 14280 -2080 15080 -2040
rect 15692 -1320 16492 -1280
rect 15692 -2040 15732 -1320
rect 16452 -2040 16492 -1320
rect 15692 -2080 16492 -2040
rect 17104 -1320 17904 -1280
rect 17104 -2040 17144 -1320
rect 17864 -2040 17904 -1320
rect 17104 -2080 17904 -2040
rect 18516 -1320 19316 -1280
rect 18516 -2040 18556 -1320
rect 19276 -2040 19316 -1320
rect 18516 -2080 19316 -2040
rect 19928 -1320 20728 -1280
rect 19928 -2040 19968 -1320
rect 20688 -2040 20728 -1320
rect 19928 -2080 20728 -2040
rect 21340 -1320 22140 -1280
rect 21340 -2040 21380 -1320
rect 22100 -2040 22140 -1320
rect 21340 -2080 22140 -2040
rect 22752 -1320 23552 -1280
rect 22752 -2040 22792 -1320
rect 23512 -2040 23552 -1320
rect 22752 -2080 23552 -2040
rect -23844 -2440 -23044 -2400
rect -23844 -3160 -23804 -2440
rect -23084 -3160 -23044 -2440
rect -23844 -3200 -23044 -3160
rect -22432 -2440 -21632 -2400
rect -22432 -3160 -22392 -2440
rect -21672 -3160 -21632 -2440
rect -22432 -3200 -21632 -3160
rect -21020 -2440 -20220 -2400
rect -21020 -3160 -20980 -2440
rect -20260 -3160 -20220 -2440
rect -21020 -3200 -20220 -3160
rect -19608 -2440 -18808 -2400
rect -19608 -3160 -19568 -2440
rect -18848 -3160 -18808 -2440
rect -19608 -3200 -18808 -3160
rect -18196 -2440 -17396 -2400
rect -18196 -3160 -18156 -2440
rect -17436 -3160 -17396 -2440
rect -18196 -3200 -17396 -3160
rect -16784 -2440 -15984 -2400
rect -16784 -3160 -16744 -2440
rect -16024 -3160 -15984 -2440
rect -16784 -3200 -15984 -3160
rect -15372 -2440 -14572 -2400
rect -15372 -3160 -15332 -2440
rect -14612 -3160 -14572 -2440
rect -15372 -3200 -14572 -3160
rect -13960 -2440 -13160 -2400
rect -13960 -3160 -13920 -2440
rect -13200 -3160 -13160 -2440
rect -13960 -3200 -13160 -3160
rect -12548 -2440 -11748 -2400
rect -12548 -3160 -12508 -2440
rect -11788 -3160 -11748 -2440
rect -12548 -3200 -11748 -3160
rect -11136 -2440 -10336 -2400
rect -11136 -3160 -11096 -2440
rect -10376 -3160 -10336 -2440
rect -11136 -3200 -10336 -3160
rect -9724 -2440 -8924 -2400
rect -9724 -3160 -9684 -2440
rect -8964 -3160 -8924 -2440
rect -9724 -3200 -8924 -3160
rect -8312 -2440 -7512 -2400
rect -8312 -3160 -8272 -2440
rect -7552 -3160 -7512 -2440
rect -8312 -3200 -7512 -3160
rect -6900 -2440 -6100 -2400
rect -6900 -3160 -6860 -2440
rect -6140 -3160 -6100 -2440
rect -6900 -3200 -6100 -3160
rect -5488 -2440 -4688 -2400
rect -5488 -3160 -5448 -2440
rect -4728 -3160 -4688 -2440
rect -5488 -3200 -4688 -3160
rect -4076 -2440 -3276 -2400
rect -4076 -3160 -4036 -2440
rect -3316 -3160 -3276 -2440
rect -4076 -3200 -3276 -3160
rect -2664 -2440 -1864 -2400
rect -2664 -3160 -2624 -2440
rect -1904 -3160 -1864 -2440
rect -2664 -3200 -1864 -3160
rect -1252 -2440 -452 -2400
rect -1252 -3160 -1212 -2440
rect -492 -3160 -452 -2440
rect -1252 -3200 -452 -3160
rect 160 -2440 960 -2400
rect 160 -3160 200 -2440
rect 920 -3160 960 -2440
rect 160 -3200 960 -3160
rect 1572 -2440 2372 -2400
rect 1572 -3160 1612 -2440
rect 2332 -3160 2372 -2440
rect 1572 -3200 2372 -3160
rect 2984 -2440 3784 -2400
rect 2984 -3160 3024 -2440
rect 3744 -3160 3784 -2440
rect 2984 -3200 3784 -3160
rect 4396 -2440 5196 -2400
rect 4396 -3160 4436 -2440
rect 5156 -3160 5196 -2440
rect 4396 -3200 5196 -3160
rect 5808 -2440 6608 -2400
rect 5808 -3160 5848 -2440
rect 6568 -3160 6608 -2440
rect 5808 -3200 6608 -3160
rect 7220 -2440 8020 -2400
rect 7220 -3160 7260 -2440
rect 7980 -3160 8020 -2440
rect 7220 -3200 8020 -3160
rect 8632 -2440 9432 -2400
rect 8632 -3160 8672 -2440
rect 9392 -3160 9432 -2440
rect 8632 -3200 9432 -3160
rect 10044 -2440 10844 -2400
rect 10044 -3160 10084 -2440
rect 10804 -3160 10844 -2440
rect 10044 -3200 10844 -3160
rect 11456 -2440 12256 -2400
rect 11456 -3160 11496 -2440
rect 12216 -3160 12256 -2440
rect 11456 -3200 12256 -3160
rect 12868 -2440 13668 -2400
rect 12868 -3160 12908 -2440
rect 13628 -3160 13668 -2440
rect 12868 -3200 13668 -3160
rect 14280 -2440 15080 -2400
rect 14280 -3160 14320 -2440
rect 15040 -3160 15080 -2440
rect 14280 -3200 15080 -3160
rect 15692 -2440 16492 -2400
rect 15692 -3160 15732 -2440
rect 16452 -3160 16492 -2440
rect 15692 -3200 16492 -3160
rect 17104 -2440 17904 -2400
rect 17104 -3160 17144 -2440
rect 17864 -3160 17904 -2440
rect 17104 -3200 17904 -3160
rect 18516 -2440 19316 -2400
rect 18516 -3160 18556 -2440
rect 19276 -3160 19316 -2440
rect 18516 -3200 19316 -3160
rect 19928 -2440 20728 -2400
rect 19928 -3160 19968 -2440
rect 20688 -3160 20728 -2440
rect 19928 -3200 20728 -3160
rect 21340 -2440 22140 -2400
rect 21340 -3160 21380 -2440
rect 22100 -3160 22140 -2440
rect 21340 -3200 22140 -3160
rect 22752 -2440 23552 -2400
rect 22752 -3160 22792 -2440
rect 23512 -3160 23552 -2440
rect 22752 -3200 23552 -3160
rect -23844 -3560 -23044 -3520
rect -23844 -4280 -23804 -3560
rect -23084 -4280 -23044 -3560
rect -23844 -4320 -23044 -4280
rect -22432 -3560 -21632 -3520
rect -22432 -4280 -22392 -3560
rect -21672 -4280 -21632 -3560
rect -22432 -4320 -21632 -4280
rect -21020 -3560 -20220 -3520
rect -21020 -4280 -20980 -3560
rect -20260 -4280 -20220 -3560
rect -21020 -4320 -20220 -4280
rect -19608 -3560 -18808 -3520
rect -19608 -4280 -19568 -3560
rect -18848 -4280 -18808 -3560
rect -19608 -4320 -18808 -4280
rect -18196 -3560 -17396 -3520
rect -18196 -4280 -18156 -3560
rect -17436 -4280 -17396 -3560
rect -18196 -4320 -17396 -4280
rect -16784 -3560 -15984 -3520
rect -16784 -4280 -16744 -3560
rect -16024 -4280 -15984 -3560
rect -16784 -4320 -15984 -4280
rect -15372 -3560 -14572 -3520
rect -15372 -4280 -15332 -3560
rect -14612 -4280 -14572 -3560
rect -15372 -4320 -14572 -4280
rect -13960 -3560 -13160 -3520
rect -13960 -4280 -13920 -3560
rect -13200 -4280 -13160 -3560
rect -13960 -4320 -13160 -4280
rect -12548 -3560 -11748 -3520
rect -12548 -4280 -12508 -3560
rect -11788 -4280 -11748 -3560
rect -12548 -4320 -11748 -4280
rect -11136 -3560 -10336 -3520
rect -11136 -4280 -11096 -3560
rect -10376 -4280 -10336 -3560
rect -11136 -4320 -10336 -4280
rect -9724 -3560 -8924 -3520
rect -9724 -4280 -9684 -3560
rect -8964 -4280 -8924 -3560
rect -9724 -4320 -8924 -4280
rect -8312 -3560 -7512 -3520
rect -8312 -4280 -8272 -3560
rect -7552 -4280 -7512 -3560
rect -8312 -4320 -7512 -4280
rect -6900 -3560 -6100 -3520
rect -6900 -4280 -6860 -3560
rect -6140 -4280 -6100 -3560
rect -6900 -4320 -6100 -4280
rect -5488 -3560 -4688 -3520
rect -5488 -4280 -5448 -3560
rect -4728 -4280 -4688 -3560
rect -5488 -4320 -4688 -4280
rect -4076 -3560 -3276 -3520
rect -4076 -4280 -4036 -3560
rect -3316 -4280 -3276 -3560
rect -4076 -4320 -3276 -4280
rect -2664 -3560 -1864 -3520
rect -2664 -4280 -2624 -3560
rect -1904 -4280 -1864 -3560
rect -2664 -4320 -1864 -4280
rect -1252 -3560 -452 -3520
rect -1252 -4280 -1212 -3560
rect -492 -4280 -452 -3560
rect -1252 -4320 -452 -4280
rect 160 -3560 960 -3520
rect 160 -4280 200 -3560
rect 920 -4280 960 -3560
rect 160 -4320 960 -4280
rect 1572 -3560 2372 -3520
rect 1572 -4280 1612 -3560
rect 2332 -4280 2372 -3560
rect 1572 -4320 2372 -4280
rect 2984 -3560 3784 -3520
rect 2984 -4280 3024 -3560
rect 3744 -4280 3784 -3560
rect 2984 -4320 3784 -4280
rect 4396 -3560 5196 -3520
rect 4396 -4280 4436 -3560
rect 5156 -4280 5196 -3560
rect 4396 -4320 5196 -4280
rect 5808 -3560 6608 -3520
rect 5808 -4280 5848 -3560
rect 6568 -4280 6608 -3560
rect 5808 -4320 6608 -4280
rect 7220 -3560 8020 -3520
rect 7220 -4280 7260 -3560
rect 7980 -4280 8020 -3560
rect 7220 -4320 8020 -4280
rect 8632 -3560 9432 -3520
rect 8632 -4280 8672 -3560
rect 9392 -4280 9432 -3560
rect 8632 -4320 9432 -4280
rect 10044 -3560 10844 -3520
rect 10044 -4280 10084 -3560
rect 10804 -4280 10844 -3560
rect 10044 -4320 10844 -4280
rect 11456 -3560 12256 -3520
rect 11456 -4280 11496 -3560
rect 12216 -4280 12256 -3560
rect 11456 -4320 12256 -4280
rect 12868 -3560 13668 -3520
rect 12868 -4280 12908 -3560
rect 13628 -4280 13668 -3560
rect 12868 -4320 13668 -4280
rect 14280 -3560 15080 -3520
rect 14280 -4280 14320 -3560
rect 15040 -4280 15080 -3560
rect 14280 -4320 15080 -4280
rect 15692 -3560 16492 -3520
rect 15692 -4280 15732 -3560
rect 16452 -4280 16492 -3560
rect 15692 -4320 16492 -4280
rect 17104 -3560 17904 -3520
rect 17104 -4280 17144 -3560
rect 17864 -4280 17904 -3560
rect 17104 -4320 17904 -4280
rect 18516 -3560 19316 -3520
rect 18516 -4280 18556 -3560
rect 19276 -4280 19316 -3560
rect 18516 -4320 19316 -4280
rect 19928 -3560 20728 -3520
rect 19928 -4280 19968 -3560
rect 20688 -4280 20728 -3560
rect 19928 -4320 20728 -4280
rect 21340 -3560 22140 -3520
rect 21340 -4280 21380 -3560
rect 22100 -4280 22140 -3560
rect 21340 -4320 22140 -4280
rect 22752 -3560 23552 -3520
rect 22752 -4280 22792 -3560
rect 23512 -4280 23552 -3560
rect 22752 -4320 23552 -4280
rect -23844 -4680 -23044 -4640
rect -23844 -5400 -23804 -4680
rect -23084 -5400 -23044 -4680
rect -23844 -5440 -23044 -5400
rect -22432 -4680 -21632 -4640
rect -22432 -5400 -22392 -4680
rect -21672 -5400 -21632 -4680
rect -22432 -5440 -21632 -5400
rect -21020 -4680 -20220 -4640
rect -21020 -5400 -20980 -4680
rect -20260 -5400 -20220 -4680
rect -21020 -5440 -20220 -5400
rect -19608 -4680 -18808 -4640
rect -19608 -5400 -19568 -4680
rect -18848 -5400 -18808 -4680
rect -19608 -5440 -18808 -5400
rect -18196 -4680 -17396 -4640
rect -18196 -5400 -18156 -4680
rect -17436 -5400 -17396 -4680
rect -18196 -5440 -17396 -5400
rect -16784 -4680 -15984 -4640
rect -16784 -5400 -16744 -4680
rect -16024 -5400 -15984 -4680
rect -16784 -5440 -15984 -5400
rect -15372 -4680 -14572 -4640
rect -15372 -5400 -15332 -4680
rect -14612 -5400 -14572 -4680
rect -15372 -5440 -14572 -5400
rect -13960 -4680 -13160 -4640
rect -13960 -5400 -13920 -4680
rect -13200 -5400 -13160 -4680
rect -13960 -5440 -13160 -5400
rect -12548 -4680 -11748 -4640
rect -12548 -5400 -12508 -4680
rect -11788 -5400 -11748 -4680
rect -12548 -5440 -11748 -5400
rect -11136 -4680 -10336 -4640
rect -11136 -5400 -11096 -4680
rect -10376 -5400 -10336 -4680
rect -11136 -5440 -10336 -5400
rect -9724 -4680 -8924 -4640
rect -9724 -5400 -9684 -4680
rect -8964 -5400 -8924 -4680
rect -9724 -5440 -8924 -5400
rect -8312 -4680 -7512 -4640
rect -8312 -5400 -8272 -4680
rect -7552 -5400 -7512 -4680
rect -8312 -5440 -7512 -5400
rect -6900 -4680 -6100 -4640
rect -6900 -5400 -6860 -4680
rect -6140 -5400 -6100 -4680
rect -6900 -5440 -6100 -5400
rect -5488 -4680 -4688 -4640
rect -5488 -5400 -5448 -4680
rect -4728 -5400 -4688 -4680
rect -5488 -5440 -4688 -5400
rect -4076 -4680 -3276 -4640
rect -4076 -5400 -4036 -4680
rect -3316 -5400 -3276 -4680
rect -4076 -5440 -3276 -5400
rect -2664 -4680 -1864 -4640
rect -2664 -5400 -2624 -4680
rect -1904 -5400 -1864 -4680
rect -2664 -5440 -1864 -5400
rect -1252 -4680 -452 -4640
rect -1252 -5400 -1212 -4680
rect -492 -5400 -452 -4680
rect -1252 -5440 -452 -5400
rect 160 -4680 960 -4640
rect 160 -5400 200 -4680
rect 920 -5400 960 -4680
rect 160 -5440 960 -5400
rect 1572 -4680 2372 -4640
rect 1572 -5400 1612 -4680
rect 2332 -5400 2372 -4680
rect 1572 -5440 2372 -5400
rect 2984 -4680 3784 -4640
rect 2984 -5400 3024 -4680
rect 3744 -5400 3784 -4680
rect 2984 -5440 3784 -5400
rect 4396 -4680 5196 -4640
rect 4396 -5400 4436 -4680
rect 5156 -5400 5196 -4680
rect 4396 -5440 5196 -5400
rect 5808 -4680 6608 -4640
rect 5808 -5400 5848 -4680
rect 6568 -5400 6608 -4680
rect 5808 -5440 6608 -5400
rect 7220 -4680 8020 -4640
rect 7220 -5400 7260 -4680
rect 7980 -5400 8020 -4680
rect 7220 -5440 8020 -5400
rect 8632 -4680 9432 -4640
rect 8632 -5400 8672 -4680
rect 9392 -5400 9432 -4680
rect 8632 -5440 9432 -5400
rect 10044 -4680 10844 -4640
rect 10044 -5400 10084 -4680
rect 10804 -5400 10844 -4680
rect 10044 -5440 10844 -5400
rect 11456 -4680 12256 -4640
rect 11456 -5400 11496 -4680
rect 12216 -5400 12256 -4680
rect 11456 -5440 12256 -5400
rect 12868 -4680 13668 -4640
rect 12868 -5400 12908 -4680
rect 13628 -5400 13668 -4680
rect 12868 -5440 13668 -5400
rect 14280 -4680 15080 -4640
rect 14280 -5400 14320 -4680
rect 15040 -5400 15080 -4680
rect 14280 -5440 15080 -5400
rect 15692 -4680 16492 -4640
rect 15692 -5400 15732 -4680
rect 16452 -5400 16492 -4680
rect 15692 -5440 16492 -5400
rect 17104 -4680 17904 -4640
rect 17104 -5400 17144 -4680
rect 17864 -5400 17904 -4680
rect 17104 -5440 17904 -5400
rect 18516 -4680 19316 -4640
rect 18516 -5400 18556 -4680
rect 19276 -5400 19316 -4680
rect 18516 -5440 19316 -5400
rect 19928 -4680 20728 -4640
rect 19928 -5400 19968 -4680
rect 20688 -5400 20728 -4680
rect 19928 -5440 20728 -5400
rect 21340 -4680 22140 -4640
rect 21340 -5400 21380 -4680
rect 22100 -5400 22140 -4680
rect 21340 -5440 22140 -5400
rect 22752 -4680 23552 -4640
rect 22752 -5400 22792 -4680
rect 23512 -5400 23552 -4680
rect 22752 -5440 23552 -5400
rect -23844 -5800 -23044 -5760
rect -23844 -6520 -23804 -5800
rect -23084 -6520 -23044 -5800
rect -23844 -6560 -23044 -6520
rect -22432 -5800 -21632 -5760
rect -22432 -6520 -22392 -5800
rect -21672 -6520 -21632 -5800
rect -22432 -6560 -21632 -6520
rect -21020 -5800 -20220 -5760
rect -21020 -6520 -20980 -5800
rect -20260 -6520 -20220 -5800
rect -21020 -6560 -20220 -6520
rect -19608 -5800 -18808 -5760
rect -19608 -6520 -19568 -5800
rect -18848 -6520 -18808 -5800
rect -19608 -6560 -18808 -6520
rect -18196 -5800 -17396 -5760
rect -18196 -6520 -18156 -5800
rect -17436 -6520 -17396 -5800
rect -18196 -6560 -17396 -6520
rect -16784 -5800 -15984 -5760
rect -16784 -6520 -16744 -5800
rect -16024 -6520 -15984 -5800
rect -16784 -6560 -15984 -6520
rect -15372 -5800 -14572 -5760
rect -15372 -6520 -15332 -5800
rect -14612 -6520 -14572 -5800
rect -15372 -6560 -14572 -6520
rect -13960 -5800 -13160 -5760
rect -13960 -6520 -13920 -5800
rect -13200 -6520 -13160 -5800
rect -13960 -6560 -13160 -6520
rect -12548 -5800 -11748 -5760
rect -12548 -6520 -12508 -5800
rect -11788 -6520 -11748 -5800
rect -12548 -6560 -11748 -6520
rect -11136 -5800 -10336 -5760
rect -11136 -6520 -11096 -5800
rect -10376 -6520 -10336 -5800
rect -11136 -6560 -10336 -6520
rect -9724 -5800 -8924 -5760
rect -9724 -6520 -9684 -5800
rect -8964 -6520 -8924 -5800
rect -9724 -6560 -8924 -6520
rect -8312 -5800 -7512 -5760
rect -8312 -6520 -8272 -5800
rect -7552 -6520 -7512 -5800
rect -8312 -6560 -7512 -6520
rect -6900 -5800 -6100 -5760
rect -6900 -6520 -6860 -5800
rect -6140 -6520 -6100 -5800
rect -6900 -6560 -6100 -6520
rect -5488 -5800 -4688 -5760
rect -5488 -6520 -5448 -5800
rect -4728 -6520 -4688 -5800
rect -5488 -6560 -4688 -6520
rect -4076 -5800 -3276 -5760
rect -4076 -6520 -4036 -5800
rect -3316 -6520 -3276 -5800
rect -4076 -6560 -3276 -6520
rect -2664 -5800 -1864 -5760
rect -2664 -6520 -2624 -5800
rect -1904 -6520 -1864 -5800
rect -2664 -6560 -1864 -6520
rect -1252 -5800 -452 -5760
rect -1252 -6520 -1212 -5800
rect -492 -6520 -452 -5800
rect -1252 -6560 -452 -6520
rect 160 -5800 960 -5760
rect 160 -6520 200 -5800
rect 920 -6520 960 -5800
rect 160 -6560 960 -6520
rect 1572 -5800 2372 -5760
rect 1572 -6520 1612 -5800
rect 2332 -6520 2372 -5800
rect 1572 -6560 2372 -6520
rect 2984 -5800 3784 -5760
rect 2984 -6520 3024 -5800
rect 3744 -6520 3784 -5800
rect 2984 -6560 3784 -6520
rect 4396 -5800 5196 -5760
rect 4396 -6520 4436 -5800
rect 5156 -6520 5196 -5800
rect 4396 -6560 5196 -6520
rect 5808 -5800 6608 -5760
rect 5808 -6520 5848 -5800
rect 6568 -6520 6608 -5800
rect 5808 -6560 6608 -6520
rect 7220 -5800 8020 -5760
rect 7220 -6520 7260 -5800
rect 7980 -6520 8020 -5800
rect 7220 -6560 8020 -6520
rect 8632 -5800 9432 -5760
rect 8632 -6520 8672 -5800
rect 9392 -6520 9432 -5800
rect 8632 -6560 9432 -6520
rect 10044 -5800 10844 -5760
rect 10044 -6520 10084 -5800
rect 10804 -6520 10844 -5800
rect 10044 -6560 10844 -6520
rect 11456 -5800 12256 -5760
rect 11456 -6520 11496 -5800
rect 12216 -6520 12256 -5800
rect 11456 -6560 12256 -6520
rect 12868 -5800 13668 -5760
rect 12868 -6520 12908 -5800
rect 13628 -6520 13668 -5800
rect 12868 -6560 13668 -6520
rect 14280 -5800 15080 -5760
rect 14280 -6520 14320 -5800
rect 15040 -6520 15080 -5800
rect 14280 -6560 15080 -6520
rect 15692 -5800 16492 -5760
rect 15692 -6520 15732 -5800
rect 16452 -6520 16492 -5800
rect 15692 -6560 16492 -6520
rect 17104 -5800 17904 -5760
rect 17104 -6520 17144 -5800
rect 17864 -6520 17904 -5800
rect 17104 -6560 17904 -6520
rect 18516 -5800 19316 -5760
rect 18516 -6520 18556 -5800
rect 19276 -6520 19316 -5800
rect 18516 -6560 19316 -6520
rect 19928 -5800 20728 -5760
rect 19928 -6520 19968 -5800
rect 20688 -6520 20728 -5800
rect 19928 -6560 20728 -6520
rect 21340 -5800 22140 -5760
rect 21340 -6520 21380 -5800
rect 22100 -6520 22140 -5800
rect 21340 -6560 22140 -6520
rect 22752 -5800 23552 -5760
rect 22752 -6520 22792 -5800
rect 23512 -6520 23552 -5800
rect 22752 -6560 23552 -6520
rect -23844 -6920 -23044 -6880
rect -23844 -7640 -23804 -6920
rect -23084 -7640 -23044 -6920
rect -23844 -7680 -23044 -7640
rect -22432 -6920 -21632 -6880
rect -22432 -7640 -22392 -6920
rect -21672 -7640 -21632 -6920
rect -22432 -7680 -21632 -7640
rect -21020 -6920 -20220 -6880
rect -21020 -7640 -20980 -6920
rect -20260 -7640 -20220 -6920
rect -21020 -7680 -20220 -7640
rect -19608 -6920 -18808 -6880
rect -19608 -7640 -19568 -6920
rect -18848 -7640 -18808 -6920
rect -19608 -7680 -18808 -7640
rect -18196 -6920 -17396 -6880
rect -18196 -7640 -18156 -6920
rect -17436 -7640 -17396 -6920
rect -18196 -7680 -17396 -7640
rect -16784 -6920 -15984 -6880
rect -16784 -7640 -16744 -6920
rect -16024 -7640 -15984 -6920
rect -16784 -7680 -15984 -7640
rect -15372 -6920 -14572 -6880
rect -15372 -7640 -15332 -6920
rect -14612 -7640 -14572 -6920
rect -15372 -7680 -14572 -7640
rect -13960 -6920 -13160 -6880
rect -13960 -7640 -13920 -6920
rect -13200 -7640 -13160 -6920
rect -13960 -7680 -13160 -7640
rect -12548 -6920 -11748 -6880
rect -12548 -7640 -12508 -6920
rect -11788 -7640 -11748 -6920
rect -12548 -7680 -11748 -7640
rect -11136 -6920 -10336 -6880
rect -11136 -7640 -11096 -6920
rect -10376 -7640 -10336 -6920
rect -11136 -7680 -10336 -7640
rect -9724 -6920 -8924 -6880
rect -9724 -7640 -9684 -6920
rect -8964 -7640 -8924 -6920
rect -9724 -7680 -8924 -7640
rect -8312 -6920 -7512 -6880
rect -8312 -7640 -8272 -6920
rect -7552 -7640 -7512 -6920
rect -8312 -7680 -7512 -7640
rect -6900 -6920 -6100 -6880
rect -6900 -7640 -6860 -6920
rect -6140 -7640 -6100 -6920
rect -6900 -7680 -6100 -7640
rect -5488 -6920 -4688 -6880
rect -5488 -7640 -5448 -6920
rect -4728 -7640 -4688 -6920
rect -5488 -7680 -4688 -7640
rect -4076 -6920 -3276 -6880
rect -4076 -7640 -4036 -6920
rect -3316 -7640 -3276 -6920
rect -4076 -7680 -3276 -7640
rect -2664 -6920 -1864 -6880
rect -2664 -7640 -2624 -6920
rect -1904 -7640 -1864 -6920
rect -2664 -7680 -1864 -7640
rect -1252 -6920 -452 -6880
rect -1252 -7640 -1212 -6920
rect -492 -7640 -452 -6920
rect -1252 -7680 -452 -7640
rect 160 -6920 960 -6880
rect 160 -7640 200 -6920
rect 920 -7640 960 -6920
rect 160 -7680 960 -7640
rect 1572 -6920 2372 -6880
rect 1572 -7640 1612 -6920
rect 2332 -7640 2372 -6920
rect 1572 -7680 2372 -7640
rect 2984 -6920 3784 -6880
rect 2984 -7640 3024 -6920
rect 3744 -7640 3784 -6920
rect 2984 -7680 3784 -7640
rect 4396 -6920 5196 -6880
rect 4396 -7640 4436 -6920
rect 5156 -7640 5196 -6920
rect 4396 -7680 5196 -7640
rect 5808 -6920 6608 -6880
rect 5808 -7640 5848 -6920
rect 6568 -7640 6608 -6920
rect 5808 -7680 6608 -7640
rect 7220 -6920 8020 -6880
rect 7220 -7640 7260 -6920
rect 7980 -7640 8020 -6920
rect 7220 -7680 8020 -7640
rect 8632 -6920 9432 -6880
rect 8632 -7640 8672 -6920
rect 9392 -7640 9432 -6920
rect 8632 -7680 9432 -7640
rect 10044 -6920 10844 -6880
rect 10044 -7640 10084 -6920
rect 10804 -7640 10844 -6920
rect 10044 -7680 10844 -7640
rect 11456 -6920 12256 -6880
rect 11456 -7640 11496 -6920
rect 12216 -7640 12256 -6920
rect 11456 -7680 12256 -7640
rect 12868 -6920 13668 -6880
rect 12868 -7640 12908 -6920
rect 13628 -7640 13668 -6920
rect 12868 -7680 13668 -7640
rect 14280 -6920 15080 -6880
rect 14280 -7640 14320 -6920
rect 15040 -7640 15080 -6920
rect 14280 -7680 15080 -7640
rect 15692 -6920 16492 -6880
rect 15692 -7640 15732 -6920
rect 16452 -7640 16492 -6920
rect 15692 -7680 16492 -7640
rect 17104 -6920 17904 -6880
rect 17104 -7640 17144 -6920
rect 17864 -7640 17904 -6920
rect 17104 -7680 17904 -7640
rect 18516 -6920 19316 -6880
rect 18516 -7640 18556 -6920
rect 19276 -7640 19316 -6920
rect 18516 -7680 19316 -7640
rect 19928 -6920 20728 -6880
rect 19928 -7640 19968 -6920
rect 20688 -7640 20728 -6920
rect 19928 -7680 20728 -7640
rect 21340 -6920 22140 -6880
rect 21340 -7640 21380 -6920
rect 22100 -7640 22140 -6920
rect 21340 -7680 22140 -7640
rect 22752 -6920 23552 -6880
rect 22752 -7640 22792 -6920
rect 23512 -7640 23552 -6920
rect 22752 -7680 23552 -7640
rect -23844 -8040 -23044 -8000
rect -23844 -8760 -23804 -8040
rect -23084 -8760 -23044 -8040
rect -23844 -8800 -23044 -8760
rect -22432 -8040 -21632 -8000
rect -22432 -8760 -22392 -8040
rect -21672 -8760 -21632 -8040
rect -22432 -8800 -21632 -8760
rect -21020 -8040 -20220 -8000
rect -21020 -8760 -20980 -8040
rect -20260 -8760 -20220 -8040
rect -21020 -8800 -20220 -8760
rect -19608 -8040 -18808 -8000
rect -19608 -8760 -19568 -8040
rect -18848 -8760 -18808 -8040
rect -19608 -8800 -18808 -8760
rect -18196 -8040 -17396 -8000
rect -18196 -8760 -18156 -8040
rect -17436 -8760 -17396 -8040
rect -18196 -8800 -17396 -8760
rect -16784 -8040 -15984 -8000
rect -16784 -8760 -16744 -8040
rect -16024 -8760 -15984 -8040
rect -16784 -8800 -15984 -8760
rect -15372 -8040 -14572 -8000
rect -15372 -8760 -15332 -8040
rect -14612 -8760 -14572 -8040
rect -15372 -8800 -14572 -8760
rect -13960 -8040 -13160 -8000
rect -13960 -8760 -13920 -8040
rect -13200 -8760 -13160 -8040
rect -13960 -8800 -13160 -8760
rect -12548 -8040 -11748 -8000
rect -12548 -8760 -12508 -8040
rect -11788 -8760 -11748 -8040
rect -12548 -8800 -11748 -8760
rect -11136 -8040 -10336 -8000
rect -11136 -8760 -11096 -8040
rect -10376 -8760 -10336 -8040
rect -11136 -8800 -10336 -8760
rect -9724 -8040 -8924 -8000
rect -9724 -8760 -9684 -8040
rect -8964 -8760 -8924 -8040
rect -9724 -8800 -8924 -8760
rect -8312 -8040 -7512 -8000
rect -8312 -8760 -8272 -8040
rect -7552 -8760 -7512 -8040
rect -8312 -8800 -7512 -8760
rect -6900 -8040 -6100 -8000
rect -6900 -8760 -6860 -8040
rect -6140 -8760 -6100 -8040
rect -6900 -8800 -6100 -8760
rect -5488 -8040 -4688 -8000
rect -5488 -8760 -5448 -8040
rect -4728 -8760 -4688 -8040
rect -5488 -8800 -4688 -8760
rect -4076 -8040 -3276 -8000
rect -4076 -8760 -4036 -8040
rect -3316 -8760 -3276 -8040
rect -4076 -8800 -3276 -8760
rect -2664 -8040 -1864 -8000
rect -2664 -8760 -2624 -8040
rect -1904 -8760 -1864 -8040
rect -2664 -8800 -1864 -8760
rect -1252 -8040 -452 -8000
rect -1252 -8760 -1212 -8040
rect -492 -8760 -452 -8040
rect -1252 -8800 -452 -8760
rect 160 -8040 960 -8000
rect 160 -8760 200 -8040
rect 920 -8760 960 -8040
rect 160 -8800 960 -8760
rect 1572 -8040 2372 -8000
rect 1572 -8760 1612 -8040
rect 2332 -8760 2372 -8040
rect 1572 -8800 2372 -8760
rect 2984 -8040 3784 -8000
rect 2984 -8760 3024 -8040
rect 3744 -8760 3784 -8040
rect 2984 -8800 3784 -8760
rect 4396 -8040 5196 -8000
rect 4396 -8760 4436 -8040
rect 5156 -8760 5196 -8040
rect 4396 -8800 5196 -8760
rect 5808 -8040 6608 -8000
rect 5808 -8760 5848 -8040
rect 6568 -8760 6608 -8040
rect 5808 -8800 6608 -8760
rect 7220 -8040 8020 -8000
rect 7220 -8760 7260 -8040
rect 7980 -8760 8020 -8040
rect 7220 -8800 8020 -8760
rect 8632 -8040 9432 -8000
rect 8632 -8760 8672 -8040
rect 9392 -8760 9432 -8040
rect 8632 -8800 9432 -8760
rect 10044 -8040 10844 -8000
rect 10044 -8760 10084 -8040
rect 10804 -8760 10844 -8040
rect 10044 -8800 10844 -8760
rect 11456 -8040 12256 -8000
rect 11456 -8760 11496 -8040
rect 12216 -8760 12256 -8040
rect 11456 -8800 12256 -8760
rect 12868 -8040 13668 -8000
rect 12868 -8760 12908 -8040
rect 13628 -8760 13668 -8040
rect 12868 -8800 13668 -8760
rect 14280 -8040 15080 -8000
rect 14280 -8760 14320 -8040
rect 15040 -8760 15080 -8040
rect 14280 -8800 15080 -8760
rect 15692 -8040 16492 -8000
rect 15692 -8760 15732 -8040
rect 16452 -8760 16492 -8040
rect 15692 -8800 16492 -8760
rect 17104 -8040 17904 -8000
rect 17104 -8760 17144 -8040
rect 17864 -8760 17904 -8040
rect 17104 -8800 17904 -8760
rect 18516 -8040 19316 -8000
rect 18516 -8760 18556 -8040
rect 19276 -8760 19316 -8040
rect 18516 -8800 19316 -8760
rect 19928 -8040 20728 -8000
rect 19928 -8760 19968 -8040
rect 20688 -8760 20728 -8040
rect 19928 -8800 20728 -8760
rect 21340 -8040 22140 -8000
rect 21340 -8760 21380 -8040
rect 22100 -8760 22140 -8040
rect 21340 -8800 22140 -8760
rect 22752 -8040 23552 -8000
rect 22752 -8760 22792 -8040
rect 23512 -8760 23552 -8040
rect 22752 -8800 23552 -8760
rect -23844 -9160 -23044 -9120
rect -23844 -9880 -23804 -9160
rect -23084 -9880 -23044 -9160
rect -23844 -9920 -23044 -9880
rect -22432 -9160 -21632 -9120
rect -22432 -9880 -22392 -9160
rect -21672 -9880 -21632 -9160
rect -22432 -9920 -21632 -9880
rect -21020 -9160 -20220 -9120
rect -21020 -9880 -20980 -9160
rect -20260 -9880 -20220 -9160
rect -21020 -9920 -20220 -9880
rect -19608 -9160 -18808 -9120
rect -19608 -9880 -19568 -9160
rect -18848 -9880 -18808 -9160
rect -19608 -9920 -18808 -9880
rect -18196 -9160 -17396 -9120
rect -18196 -9880 -18156 -9160
rect -17436 -9880 -17396 -9160
rect -18196 -9920 -17396 -9880
rect -16784 -9160 -15984 -9120
rect -16784 -9880 -16744 -9160
rect -16024 -9880 -15984 -9160
rect -16784 -9920 -15984 -9880
rect -15372 -9160 -14572 -9120
rect -15372 -9880 -15332 -9160
rect -14612 -9880 -14572 -9160
rect -15372 -9920 -14572 -9880
rect -13960 -9160 -13160 -9120
rect -13960 -9880 -13920 -9160
rect -13200 -9880 -13160 -9160
rect -13960 -9920 -13160 -9880
rect -12548 -9160 -11748 -9120
rect -12548 -9880 -12508 -9160
rect -11788 -9880 -11748 -9160
rect -12548 -9920 -11748 -9880
rect -11136 -9160 -10336 -9120
rect -11136 -9880 -11096 -9160
rect -10376 -9880 -10336 -9160
rect -11136 -9920 -10336 -9880
rect -9724 -9160 -8924 -9120
rect -9724 -9880 -9684 -9160
rect -8964 -9880 -8924 -9160
rect -9724 -9920 -8924 -9880
rect -8312 -9160 -7512 -9120
rect -8312 -9880 -8272 -9160
rect -7552 -9880 -7512 -9160
rect -8312 -9920 -7512 -9880
rect -6900 -9160 -6100 -9120
rect -6900 -9880 -6860 -9160
rect -6140 -9880 -6100 -9160
rect -6900 -9920 -6100 -9880
rect -5488 -9160 -4688 -9120
rect -5488 -9880 -5448 -9160
rect -4728 -9880 -4688 -9160
rect -5488 -9920 -4688 -9880
rect -4076 -9160 -3276 -9120
rect -4076 -9880 -4036 -9160
rect -3316 -9880 -3276 -9160
rect -4076 -9920 -3276 -9880
rect -2664 -9160 -1864 -9120
rect -2664 -9880 -2624 -9160
rect -1904 -9880 -1864 -9160
rect -2664 -9920 -1864 -9880
rect -1252 -9160 -452 -9120
rect -1252 -9880 -1212 -9160
rect -492 -9880 -452 -9160
rect -1252 -9920 -452 -9880
rect 160 -9160 960 -9120
rect 160 -9880 200 -9160
rect 920 -9880 960 -9160
rect 160 -9920 960 -9880
rect 1572 -9160 2372 -9120
rect 1572 -9880 1612 -9160
rect 2332 -9880 2372 -9160
rect 1572 -9920 2372 -9880
rect 2984 -9160 3784 -9120
rect 2984 -9880 3024 -9160
rect 3744 -9880 3784 -9160
rect 2984 -9920 3784 -9880
rect 4396 -9160 5196 -9120
rect 4396 -9880 4436 -9160
rect 5156 -9880 5196 -9160
rect 4396 -9920 5196 -9880
rect 5808 -9160 6608 -9120
rect 5808 -9880 5848 -9160
rect 6568 -9880 6608 -9160
rect 5808 -9920 6608 -9880
rect 7220 -9160 8020 -9120
rect 7220 -9880 7260 -9160
rect 7980 -9880 8020 -9160
rect 7220 -9920 8020 -9880
rect 8632 -9160 9432 -9120
rect 8632 -9880 8672 -9160
rect 9392 -9880 9432 -9160
rect 8632 -9920 9432 -9880
rect 10044 -9160 10844 -9120
rect 10044 -9880 10084 -9160
rect 10804 -9880 10844 -9160
rect 10044 -9920 10844 -9880
rect 11456 -9160 12256 -9120
rect 11456 -9880 11496 -9160
rect 12216 -9880 12256 -9160
rect 11456 -9920 12256 -9880
rect 12868 -9160 13668 -9120
rect 12868 -9880 12908 -9160
rect 13628 -9880 13668 -9160
rect 12868 -9920 13668 -9880
rect 14280 -9160 15080 -9120
rect 14280 -9880 14320 -9160
rect 15040 -9880 15080 -9160
rect 14280 -9920 15080 -9880
rect 15692 -9160 16492 -9120
rect 15692 -9880 15732 -9160
rect 16452 -9880 16492 -9160
rect 15692 -9920 16492 -9880
rect 17104 -9160 17904 -9120
rect 17104 -9880 17144 -9160
rect 17864 -9880 17904 -9160
rect 17104 -9920 17904 -9880
rect 18516 -9160 19316 -9120
rect 18516 -9880 18556 -9160
rect 19276 -9880 19316 -9160
rect 18516 -9920 19316 -9880
rect 19928 -9160 20728 -9120
rect 19928 -9880 19968 -9160
rect 20688 -9880 20728 -9160
rect 19928 -9920 20728 -9880
rect 21340 -9160 22140 -9120
rect 21340 -9880 21380 -9160
rect 22100 -9880 22140 -9160
rect 21340 -9920 22140 -9880
rect 22752 -9160 23552 -9120
rect 22752 -9880 22792 -9160
rect 23512 -9880 23552 -9160
rect 22752 -9920 23552 -9880
rect -23844 -10280 -23044 -10240
rect -23844 -11000 -23804 -10280
rect -23084 -11000 -23044 -10280
rect -23844 -11040 -23044 -11000
rect -22432 -10280 -21632 -10240
rect -22432 -11000 -22392 -10280
rect -21672 -11000 -21632 -10280
rect -22432 -11040 -21632 -11000
rect -21020 -10280 -20220 -10240
rect -21020 -11000 -20980 -10280
rect -20260 -11000 -20220 -10280
rect -21020 -11040 -20220 -11000
rect -19608 -10280 -18808 -10240
rect -19608 -11000 -19568 -10280
rect -18848 -11000 -18808 -10280
rect -19608 -11040 -18808 -11000
rect -18196 -10280 -17396 -10240
rect -18196 -11000 -18156 -10280
rect -17436 -11000 -17396 -10280
rect -18196 -11040 -17396 -11000
rect -16784 -10280 -15984 -10240
rect -16784 -11000 -16744 -10280
rect -16024 -11000 -15984 -10280
rect -16784 -11040 -15984 -11000
rect -15372 -10280 -14572 -10240
rect -15372 -11000 -15332 -10280
rect -14612 -11000 -14572 -10280
rect -15372 -11040 -14572 -11000
rect -13960 -10280 -13160 -10240
rect -13960 -11000 -13920 -10280
rect -13200 -11000 -13160 -10280
rect -13960 -11040 -13160 -11000
rect -12548 -10280 -11748 -10240
rect -12548 -11000 -12508 -10280
rect -11788 -11000 -11748 -10280
rect -12548 -11040 -11748 -11000
rect -11136 -10280 -10336 -10240
rect -11136 -11000 -11096 -10280
rect -10376 -11000 -10336 -10280
rect -11136 -11040 -10336 -11000
rect -9724 -10280 -8924 -10240
rect -9724 -11000 -9684 -10280
rect -8964 -11000 -8924 -10280
rect -9724 -11040 -8924 -11000
rect -8312 -10280 -7512 -10240
rect -8312 -11000 -8272 -10280
rect -7552 -11000 -7512 -10280
rect -8312 -11040 -7512 -11000
rect -6900 -10280 -6100 -10240
rect -6900 -11000 -6860 -10280
rect -6140 -11000 -6100 -10280
rect -6900 -11040 -6100 -11000
rect -5488 -10280 -4688 -10240
rect -5488 -11000 -5448 -10280
rect -4728 -11000 -4688 -10280
rect -5488 -11040 -4688 -11000
rect -4076 -10280 -3276 -10240
rect -4076 -11000 -4036 -10280
rect -3316 -11000 -3276 -10280
rect -4076 -11040 -3276 -11000
rect -2664 -10280 -1864 -10240
rect -2664 -11000 -2624 -10280
rect -1904 -11000 -1864 -10280
rect -2664 -11040 -1864 -11000
rect -1252 -10280 -452 -10240
rect -1252 -11000 -1212 -10280
rect -492 -11000 -452 -10280
rect -1252 -11040 -452 -11000
rect 160 -10280 960 -10240
rect 160 -11000 200 -10280
rect 920 -11000 960 -10280
rect 160 -11040 960 -11000
rect 1572 -10280 2372 -10240
rect 1572 -11000 1612 -10280
rect 2332 -11000 2372 -10280
rect 1572 -11040 2372 -11000
rect 2984 -10280 3784 -10240
rect 2984 -11000 3024 -10280
rect 3744 -11000 3784 -10280
rect 2984 -11040 3784 -11000
rect 4396 -10280 5196 -10240
rect 4396 -11000 4436 -10280
rect 5156 -11000 5196 -10280
rect 4396 -11040 5196 -11000
rect 5808 -10280 6608 -10240
rect 5808 -11000 5848 -10280
rect 6568 -11000 6608 -10280
rect 5808 -11040 6608 -11000
rect 7220 -10280 8020 -10240
rect 7220 -11000 7260 -10280
rect 7980 -11000 8020 -10280
rect 7220 -11040 8020 -11000
rect 8632 -10280 9432 -10240
rect 8632 -11000 8672 -10280
rect 9392 -11000 9432 -10280
rect 8632 -11040 9432 -11000
rect 10044 -10280 10844 -10240
rect 10044 -11000 10084 -10280
rect 10804 -11000 10844 -10280
rect 10044 -11040 10844 -11000
rect 11456 -10280 12256 -10240
rect 11456 -11000 11496 -10280
rect 12216 -11000 12256 -10280
rect 11456 -11040 12256 -11000
rect 12868 -10280 13668 -10240
rect 12868 -11000 12908 -10280
rect 13628 -11000 13668 -10280
rect 12868 -11040 13668 -11000
rect 14280 -10280 15080 -10240
rect 14280 -11000 14320 -10280
rect 15040 -11000 15080 -10280
rect 14280 -11040 15080 -11000
rect 15692 -10280 16492 -10240
rect 15692 -11000 15732 -10280
rect 16452 -11000 16492 -10280
rect 15692 -11040 16492 -11000
rect 17104 -10280 17904 -10240
rect 17104 -11000 17144 -10280
rect 17864 -11000 17904 -10280
rect 17104 -11040 17904 -11000
rect 18516 -10280 19316 -10240
rect 18516 -11000 18556 -10280
rect 19276 -11000 19316 -10280
rect 18516 -11040 19316 -11000
rect 19928 -10280 20728 -10240
rect 19928 -11000 19968 -10280
rect 20688 -11000 20728 -10280
rect 19928 -11040 20728 -11000
rect 21340 -10280 22140 -10240
rect 21340 -11000 21380 -10280
rect 22100 -11000 22140 -10280
rect 21340 -11040 22140 -11000
rect 22752 -10280 23552 -10240
rect 22752 -11000 22792 -10280
rect 23512 -11000 23552 -10280
rect 22752 -11040 23552 -11000
rect -23844 -11400 -23044 -11360
rect -23844 -12120 -23804 -11400
rect -23084 -12120 -23044 -11400
rect -23844 -12160 -23044 -12120
rect -22432 -11400 -21632 -11360
rect -22432 -12120 -22392 -11400
rect -21672 -12120 -21632 -11400
rect -22432 -12160 -21632 -12120
rect -21020 -11400 -20220 -11360
rect -21020 -12120 -20980 -11400
rect -20260 -12120 -20220 -11400
rect -21020 -12160 -20220 -12120
rect -19608 -11400 -18808 -11360
rect -19608 -12120 -19568 -11400
rect -18848 -12120 -18808 -11400
rect -19608 -12160 -18808 -12120
rect -18196 -11400 -17396 -11360
rect -18196 -12120 -18156 -11400
rect -17436 -12120 -17396 -11400
rect -18196 -12160 -17396 -12120
rect -16784 -11400 -15984 -11360
rect -16784 -12120 -16744 -11400
rect -16024 -12120 -15984 -11400
rect -16784 -12160 -15984 -12120
rect -15372 -11400 -14572 -11360
rect -15372 -12120 -15332 -11400
rect -14612 -12120 -14572 -11400
rect -15372 -12160 -14572 -12120
rect -13960 -11400 -13160 -11360
rect -13960 -12120 -13920 -11400
rect -13200 -12120 -13160 -11400
rect -13960 -12160 -13160 -12120
rect -12548 -11400 -11748 -11360
rect -12548 -12120 -12508 -11400
rect -11788 -12120 -11748 -11400
rect -12548 -12160 -11748 -12120
rect -11136 -11400 -10336 -11360
rect -11136 -12120 -11096 -11400
rect -10376 -12120 -10336 -11400
rect -11136 -12160 -10336 -12120
rect -9724 -11400 -8924 -11360
rect -9724 -12120 -9684 -11400
rect -8964 -12120 -8924 -11400
rect -9724 -12160 -8924 -12120
rect -8312 -11400 -7512 -11360
rect -8312 -12120 -8272 -11400
rect -7552 -12120 -7512 -11400
rect -8312 -12160 -7512 -12120
rect -6900 -11400 -6100 -11360
rect -6900 -12120 -6860 -11400
rect -6140 -12120 -6100 -11400
rect -6900 -12160 -6100 -12120
rect -5488 -11400 -4688 -11360
rect -5488 -12120 -5448 -11400
rect -4728 -12120 -4688 -11400
rect -5488 -12160 -4688 -12120
rect -4076 -11400 -3276 -11360
rect -4076 -12120 -4036 -11400
rect -3316 -12120 -3276 -11400
rect -4076 -12160 -3276 -12120
rect -2664 -11400 -1864 -11360
rect -2664 -12120 -2624 -11400
rect -1904 -12120 -1864 -11400
rect -2664 -12160 -1864 -12120
rect -1252 -11400 -452 -11360
rect -1252 -12120 -1212 -11400
rect -492 -12120 -452 -11400
rect -1252 -12160 -452 -12120
rect 160 -11400 960 -11360
rect 160 -12120 200 -11400
rect 920 -12120 960 -11400
rect 160 -12160 960 -12120
rect 1572 -11400 2372 -11360
rect 1572 -12120 1612 -11400
rect 2332 -12120 2372 -11400
rect 1572 -12160 2372 -12120
rect 2984 -11400 3784 -11360
rect 2984 -12120 3024 -11400
rect 3744 -12120 3784 -11400
rect 2984 -12160 3784 -12120
rect 4396 -11400 5196 -11360
rect 4396 -12120 4436 -11400
rect 5156 -12120 5196 -11400
rect 4396 -12160 5196 -12120
rect 5808 -11400 6608 -11360
rect 5808 -12120 5848 -11400
rect 6568 -12120 6608 -11400
rect 5808 -12160 6608 -12120
rect 7220 -11400 8020 -11360
rect 7220 -12120 7260 -11400
rect 7980 -12120 8020 -11400
rect 7220 -12160 8020 -12120
rect 8632 -11400 9432 -11360
rect 8632 -12120 8672 -11400
rect 9392 -12120 9432 -11400
rect 8632 -12160 9432 -12120
rect 10044 -11400 10844 -11360
rect 10044 -12120 10084 -11400
rect 10804 -12120 10844 -11400
rect 10044 -12160 10844 -12120
rect 11456 -11400 12256 -11360
rect 11456 -12120 11496 -11400
rect 12216 -12120 12256 -11400
rect 11456 -12160 12256 -12120
rect 12868 -11400 13668 -11360
rect 12868 -12120 12908 -11400
rect 13628 -12120 13668 -11400
rect 12868 -12160 13668 -12120
rect 14280 -11400 15080 -11360
rect 14280 -12120 14320 -11400
rect 15040 -12120 15080 -11400
rect 14280 -12160 15080 -12120
rect 15692 -11400 16492 -11360
rect 15692 -12120 15732 -11400
rect 16452 -12120 16492 -11400
rect 15692 -12160 16492 -12120
rect 17104 -11400 17904 -11360
rect 17104 -12120 17144 -11400
rect 17864 -12120 17904 -11400
rect 17104 -12160 17904 -12120
rect 18516 -11400 19316 -11360
rect 18516 -12120 18556 -11400
rect 19276 -12120 19316 -11400
rect 18516 -12160 19316 -12120
rect 19928 -11400 20728 -11360
rect 19928 -12120 19968 -11400
rect 20688 -12120 20728 -11400
rect 19928 -12160 20728 -12120
rect 21340 -11400 22140 -11360
rect 21340 -12120 21380 -11400
rect 22100 -12120 22140 -11400
rect 21340 -12160 22140 -12120
rect 22752 -11400 23552 -11360
rect 22752 -12120 22792 -11400
rect 23512 -12120 23552 -11400
rect 22752 -12160 23552 -12120
rect -23844 -12520 -23044 -12480
rect -23844 -13240 -23804 -12520
rect -23084 -13240 -23044 -12520
rect -23844 -13280 -23044 -13240
rect -22432 -12520 -21632 -12480
rect -22432 -13240 -22392 -12520
rect -21672 -13240 -21632 -12520
rect -22432 -13280 -21632 -13240
rect -21020 -12520 -20220 -12480
rect -21020 -13240 -20980 -12520
rect -20260 -13240 -20220 -12520
rect -21020 -13280 -20220 -13240
rect -19608 -12520 -18808 -12480
rect -19608 -13240 -19568 -12520
rect -18848 -13240 -18808 -12520
rect -19608 -13280 -18808 -13240
rect -18196 -12520 -17396 -12480
rect -18196 -13240 -18156 -12520
rect -17436 -13240 -17396 -12520
rect -18196 -13280 -17396 -13240
rect -16784 -12520 -15984 -12480
rect -16784 -13240 -16744 -12520
rect -16024 -13240 -15984 -12520
rect -16784 -13280 -15984 -13240
rect -15372 -12520 -14572 -12480
rect -15372 -13240 -15332 -12520
rect -14612 -13240 -14572 -12520
rect -15372 -13280 -14572 -13240
rect -13960 -12520 -13160 -12480
rect -13960 -13240 -13920 -12520
rect -13200 -13240 -13160 -12520
rect -13960 -13280 -13160 -13240
rect -12548 -12520 -11748 -12480
rect -12548 -13240 -12508 -12520
rect -11788 -13240 -11748 -12520
rect -12548 -13280 -11748 -13240
rect -11136 -12520 -10336 -12480
rect -11136 -13240 -11096 -12520
rect -10376 -13240 -10336 -12520
rect -11136 -13280 -10336 -13240
rect -9724 -12520 -8924 -12480
rect -9724 -13240 -9684 -12520
rect -8964 -13240 -8924 -12520
rect -9724 -13280 -8924 -13240
rect -8312 -12520 -7512 -12480
rect -8312 -13240 -8272 -12520
rect -7552 -13240 -7512 -12520
rect -8312 -13280 -7512 -13240
rect -6900 -12520 -6100 -12480
rect -6900 -13240 -6860 -12520
rect -6140 -13240 -6100 -12520
rect -6900 -13280 -6100 -13240
rect -5488 -12520 -4688 -12480
rect -5488 -13240 -5448 -12520
rect -4728 -13240 -4688 -12520
rect -5488 -13280 -4688 -13240
rect -4076 -12520 -3276 -12480
rect -4076 -13240 -4036 -12520
rect -3316 -13240 -3276 -12520
rect -4076 -13280 -3276 -13240
rect -2664 -12520 -1864 -12480
rect -2664 -13240 -2624 -12520
rect -1904 -13240 -1864 -12520
rect -2664 -13280 -1864 -13240
rect -1252 -12520 -452 -12480
rect -1252 -13240 -1212 -12520
rect -492 -13240 -452 -12520
rect -1252 -13280 -452 -13240
rect 160 -12520 960 -12480
rect 160 -13240 200 -12520
rect 920 -13240 960 -12520
rect 160 -13280 960 -13240
rect 1572 -12520 2372 -12480
rect 1572 -13240 1612 -12520
rect 2332 -13240 2372 -12520
rect 1572 -13280 2372 -13240
rect 2984 -12520 3784 -12480
rect 2984 -13240 3024 -12520
rect 3744 -13240 3784 -12520
rect 2984 -13280 3784 -13240
rect 4396 -12520 5196 -12480
rect 4396 -13240 4436 -12520
rect 5156 -13240 5196 -12520
rect 4396 -13280 5196 -13240
rect 5808 -12520 6608 -12480
rect 5808 -13240 5848 -12520
rect 6568 -13240 6608 -12520
rect 5808 -13280 6608 -13240
rect 7220 -12520 8020 -12480
rect 7220 -13240 7260 -12520
rect 7980 -13240 8020 -12520
rect 7220 -13280 8020 -13240
rect 8632 -12520 9432 -12480
rect 8632 -13240 8672 -12520
rect 9392 -13240 9432 -12520
rect 8632 -13280 9432 -13240
rect 10044 -12520 10844 -12480
rect 10044 -13240 10084 -12520
rect 10804 -13240 10844 -12520
rect 10044 -13280 10844 -13240
rect 11456 -12520 12256 -12480
rect 11456 -13240 11496 -12520
rect 12216 -13240 12256 -12520
rect 11456 -13280 12256 -13240
rect 12868 -12520 13668 -12480
rect 12868 -13240 12908 -12520
rect 13628 -13240 13668 -12520
rect 12868 -13280 13668 -13240
rect 14280 -12520 15080 -12480
rect 14280 -13240 14320 -12520
rect 15040 -13240 15080 -12520
rect 14280 -13280 15080 -13240
rect 15692 -12520 16492 -12480
rect 15692 -13240 15732 -12520
rect 16452 -13240 16492 -12520
rect 15692 -13280 16492 -13240
rect 17104 -12520 17904 -12480
rect 17104 -13240 17144 -12520
rect 17864 -13240 17904 -12520
rect 17104 -13280 17904 -13240
rect 18516 -12520 19316 -12480
rect 18516 -13240 18556 -12520
rect 19276 -13240 19316 -12520
rect 18516 -13280 19316 -13240
rect 19928 -12520 20728 -12480
rect 19928 -13240 19968 -12520
rect 20688 -13240 20728 -12520
rect 19928 -13280 20728 -13240
rect 21340 -12520 22140 -12480
rect 21340 -13240 21380 -12520
rect 22100 -13240 22140 -12520
rect 21340 -13280 22140 -13240
rect 22752 -12520 23552 -12480
rect 22752 -13240 22792 -12520
rect 23512 -13240 23552 -12520
rect 22752 -13280 23552 -13240
rect -23844 -13640 -23044 -13600
rect -23844 -14360 -23804 -13640
rect -23084 -14360 -23044 -13640
rect -23844 -14400 -23044 -14360
rect -22432 -13640 -21632 -13600
rect -22432 -14360 -22392 -13640
rect -21672 -14360 -21632 -13640
rect -22432 -14400 -21632 -14360
rect -21020 -13640 -20220 -13600
rect -21020 -14360 -20980 -13640
rect -20260 -14360 -20220 -13640
rect -21020 -14400 -20220 -14360
rect -19608 -13640 -18808 -13600
rect -19608 -14360 -19568 -13640
rect -18848 -14360 -18808 -13640
rect -19608 -14400 -18808 -14360
rect -18196 -13640 -17396 -13600
rect -18196 -14360 -18156 -13640
rect -17436 -14360 -17396 -13640
rect -18196 -14400 -17396 -14360
rect -16784 -13640 -15984 -13600
rect -16784 -14360 -16744 -13640
rect -16024 -14360 -15984 -13640
rect -16784 -14400 -15984 -14360
rect -15372 -13640 -14572 -13600
rect -15372 -14360 -15332 -13640
rect -14612 -14360 -14572 -13640
rect -15372 -14400 -14572 -14360
rect -13960 -13640 -13160 -13600
rect -13960 -14360 -13920 -13640
rect -13200 -14360 -13160 -13640
rect -13960 -14400 -13160 -14360
rect -12548 -13640 -11748 -13600
rect -12548 -14360 -12508 -13640
rect -11788 -14360 -11748 -13640
rect -12548 -14400 -11748 -14360
rect -11136 -13640 -10336 -13600
rect -11136 -14360 -11096 -13640
rect -10376 -14360 -10336 -13640
rect -11136 -14400 -10336 -14360
rect -9724 -13640 -8924 -13600
rect -9724 -14360 -9684 -13640
rect -8964 -14360 -8924 -13640
rect -9724 -14400 -8924 -14360
rect -8312 -13640 -7512 -13600
rect -8312 -14360 -8272 -13640
rect -7552 -14360 -7512 -13640
rect -8312 -14400 -7512 -14360
rect -6900 -13640 -6100 -13600
rect -6900 -14360 -6860 -13640
rect -6140 -14360 -6100 -13640
rect -6900 -14400 -6100 -14360
rect -5488 -13640 -4688 -13600
rect -5488 -14360 -5448 -13640
rect -4728 -14360 -4688 -13640
rect -5488 -14400 -4688 -14360
rect -4076 -13640 -3276 -13600
rect -4076 -14360 -4036 -13640
rect -3316 -14360 -3276 -13640
rect -4076 -14400 -3276 -14360
rect -2664 -13640 -1864 -13600
rect -2664 -14360 -2624 -13640
rect -1904 -14360 -1864 -13640
rect -2664 -14400 -1864 -14360
rect -1252 -13640 -452 -13600
rect -1252 -14360 -1212 -13640
rect -492 -14360 -452 -13640
rect -1252 -14400 -452 -14360
rect 160 -13640 960 -13600
rect 160 -14360 200 -13640
rect 920 -14360 960 -13640
rect 160 -14400 960 -14360
rect 1572 -13640 2372 -13600
rect 1572 -14360 1612 -13640
rect 2332 -14360 2372 -13640
rect 1572 -14400 2372 -14360
rect 2984 -13640 3784 -13600
rect 2984 -14360 3024 -13640
rect 3744 -14360 3784 -13640
rect 2984 -14400 3784 -14360
rect 4396 -13640 5196 -13600
rect 4396 -14360 4436 -13640
rect 5156 -14360 5196 -13640
rect 4396 -14400 5196 -14360
rect 5808 -13640 6608 -13600
rect 5808 -14360 5848 -13640
rect 6568 -14360 6608 -13640
rect 5808 -14400 6608 -14360
rect 7220 -13640 8020 -13600
rect 7220 -14360 7260 -13640
rect 7980 -14360 8020 -13640
rect 7220 -14400 8020 -14360
rect 8632 -13640 9432 -13600
rect 8632 -14360 8672 -13640
rect 9392 -14360 9432 -13640
rect 8632 -14400 9432 -14360
rect 10044 -13640 10844 -13600
rect 10044 -14360 10084 -13640
rect 10804 -14360 10844 -13640
rect 10044 -14400 10844 -14360
rect 11456 -13640 12256 -13600
rect 11456 -14360 11496 -13640
rect 12216 -14360 12256 -13640
rect 11456 -14400 12256 -14360
rect 12868 -13640 13668 -13600
rect 12868 -14360 12908 -13640
rect 13628 -14360 13668 -13640
rect 12868 -14400 13668 -14360
rect 14280 -13640 15080 -13600
rect 14280 -14360 14320 -13640
rect 15040 -14360 15080 -13640
rect 14280 -14400 15080 -14360
rect 15692 -13640 16492 -13600
rect 15692 -14360 15732 -13640
rect 16452 -14360 16492 -13640
rect 15692 -14400 16492 -14360
rect 17104 -13640 17904 -13600
rect 17104 -14360 17144 -13640
rect 17864 -14360 17904 -13640
rect 17104 -14400 17904 -14360
rect 18516 -13640 19316 -13600
rect 18516 -14360 18556 -13640
rect 19276 -14360 19316 -13640
rect 18516 -14400 19316 -14360
rect 19928 -13640 20728 -13600
rect 19928 -14360 19968 -13640
rect 20688 -14360 20728 -13640
rect 19928 -14400 20728 -14360
rect 21340 -13640 22140 -13600
rect 21340 -14360 21380 -13640
rect 22100 -14360 22140 -13640
rect 21340 -14400 22140 -14360
rect 22752 -13640 23552 -13600
rect 22752 -14360 22792 -13640
rect 23512 -14360 23552 -13640
rect 22752 -14400 23552 -14360
rect -23844 -14760 -23044 -14720
rect -23844 -15480 -23804 -14760
rect -23084 -15480 -23044 -14760
rect -23844 -15520 -23044 -15480
rect -22432 -14760 -21632 -14720
rect -22432 -15480 -22392 -14760
rect -21672 -15480 -21632 -14760
rect -22432 -15520 -21632 -15480
rect -21020 -14760 -20220 -14720
rect -21020 -15480 -20980 -14760
rect -20260 -15480 -20220 -14760
rect -21020 -15520 -20220 -15480
rect -19608 -14760 -18808 -14720
rect -19608 -15480 -19568 -14760
rect -18848 -15480 -18808 -14760
rect -19608 -15520 -18808 -15480
rect -18196 -14760 -17396 -14720
rect -18196 -15480 -18156 -14760
rect -17436 -15480 -17396 -14760
rect -18196 -15520 -17396 -15480
rect -16784 -14760 -15984 -14720
rect -16784 -15480 -16744 -14760
rect -16024 -15480 -15984 -14760
rect -16784 -15520 -15984 -15480
rect -15372 -14760 -14572 -14720
rect -15372 -15480 -15332 -14760
rect -14612 -15480 -14572 -14760
rect -15372 -15520 -14572 -15480
rect -13960 -14760 -13160 -14720
rect -13960 -15480 -13920 -14760
rect -13200 -15480 -13160 -14760
rect -13960 -15520 -13160 -15480
rect -12548 -14760 -11748 -14720
rect -12548 -15480 -12508 -14760
rect -11788 -15480 -11748 -14760
rect -12548 -15520 -11748 -15480
rect -11136 -14760 -10336 -14720
rect -11136 -15480 -11096 -14760
rect -10376 -15480 -10336 -14760
rect -11136 -15520 -10336 -15480
rect -9724 -14760 -8924 -14720
rect -9724 -15480 -9684 -14760
rect -8964 -15480 -8924 -14760
rect -9724 -15520 -8924 -15480
rect -8312 -14760 -7512 -14720
rect -8312 -15480 -8272 -14760
rect -7552 -15480 -7512 -14760
rect -8312 -15520 -7512 -15480
rect -6900 -14760 -6100 -14720
rect -6900 -15480 -6860 -14760
rect -6140 -15480 -6100 -14760
rect -6900 -15520 -6100 -15480
rect -5488 -14760 -4688 -14720
rect -5488 -15480 -5448 -14760
rect -4728 -15480 -4688 -14760
rect -5488 -15520 -4688 -15480
rect -4076 -14760 -3276 -14720
rect -4076 -15480 -4036 -14760
rect -3316 -15480 -3276 -14760
rect -4076 -15520 -3276 -15480
rect -2664 -14760 -1864 -14720
rect -2664 -15480 -2624 -14760
rect -1904 -15480 -1864 -14760
rect -2664 -15520 -1864 -15480
rect -1252 -14760 -452 -14720
rect -1252 -15480 -1212 -14760
rect -492 -15480 -452 -14760
rect -1252 -15520 -452 -15480
rect 160 -14760 960 -14720
rect 160 -15480 200 -14760
rect 920 -15480 960 -14760
rect 160 -15520 960 -15480
rect 1572 -14760 2372 -14720
rect 1572 -15480 1612 -14760
rect 2332 -15480 2372 -14760
rect 1572 -15520 2372 -15480
rect 2984 -14760 3784 -14720
rect 2984 -15480 3024 -14760
rect 3744 -15480 3784 -14760
rect 2984 -15520 3784 -15480
rect 4396 -14760 5196 -14720
rect 4396 -15480 4436 -14760
rect 5156 -15480 5196 -14760
rect 4396 -15520 5196 -15480
rect 5808 -14760 6608 -14720
rect 5808 -15480 5848 -14760
rect 6568 -15480 6608 -14760
rect 5808 -15520 6608 -15480
rect 7220 -14760 8020 -14720
rect 7220 -15480 7260 -14760
rect 7980 -15480 8020 -14760
rect 7220 -15520 8020 -15480
rect 8632 -14760 9432 -14720
rect 8632 -15480 8672 -14760
rect 9392 -15480 9432 -14760
rect 8632 -15520 9432 -15480
rect 10044 -14760 10844 -14720
rect 10044 -15480 10084 -14760
rect 10804 -15480 10844 -14760
rect 10044 -15520 10844 -15480
rect 11456 -14760 12256 -14720
rect 11456 -15480 11496 -14760
rect 12216 -15480 12256 -14760
rect 11456 -15520 12256 -15480
rect 12868 -14760 13668 -14720
rect 12868 -15480 12908 -14760
rect 13628 -15480 13668 -14760
rect 12868 -15520 13668 -15480
rect 14280 -14760 15080 -14720
rect 14280 -15480 14320 -14760
rect 15040 -15480 15080 -14760
rect 14280 -15520 15080 -15480
rect 15692 -14760 16492 -14720
rect 15692 -15480 15732 -14760
rect 16452 -15480 16492 -14760
rect 15692 -15520 16492 -15480
rect 17104 -14760 17904 -14720
rect 17104 -15480 17144 -14760
rect 17864 -15480 17904 -14760
rect 17104 -15520 17904 -15480
rect 18516 -14760 19316 -14720
rect 18516 -15480 18556 -14760
rect 19276 -15480 19316 -14760
rect 18516 -15520 19316 -15480
rect 19928 -14760 20728 -14720
rect 19928 -15480 19968 -14760
rect 20688 -15480 20728 -14760
rect 19928 -15520 20728 -15480
rect 21340 -14760 22140 -14720
rect 21340 -15480 21380 -14760
rect 22100 -15480 22140 -14760
rect 21340 -15520 22140 -15480
rect 22752 -14760 23552 -14720
rect 22752 -15480 22792 -14760
rect 23512 -15480 23552 -14760
rect 22752 -15520 23552 -15480
rect -23844 -15880 -23044 -15840
rect -23844 -16600 -23804 -15880
rect -23084 -16600 -23044 -15880
rect -23844 -16640 -23044 -16600
rect -22432 -15880 -21632 -15840
rect -22432 -16600 -22392 -15880
rect -21672 -16600 -21632 -15880
rect -22432 -16640 -21632 -16600
rect -21020 -15880 -20220 -15840
rect -21020 -16600 -20980 -15880
rect -20260 -16600 -20220 -15880
rect -21020 -16640 -20220 -16600
rect -19608 -15880 -18808 -15840
rect -19608 -16600 -19568 -15880
rect -18848 -16600 -18808 -15880
rect -19608 -16640 -18808 -16600
rect -18196 -15880 -17396 -15840
rect -18196 -16600 -18156 -15880
rect -17436 -16600 -17396 -15880
rect -18196 -16640 -17396 -16600
rect -16784 -15880 -15984 -15840
rect -16784 -16600 -16744 -15880
rect -16024 -16600 -15984 -15880
rect -16784 -16640 -15984 -16600
rect -15372 -15880 -14572 -15840
rect -15372 -16600 -15332 -15880
rect -14612 -16600 -14572 -15880
rect -15372 -16640 -14572 -16600
rect -13960 -15880 -13160 -15840
rect -13960 -16600 -13920 -15880
rect -13200 -16600 -13160 -15880
rect -13960 -16640 -13160 -16600
rect -12548 -15880 -11748 -15840
rect -12548 -16600 -12508 -15880
rect -11788 -16600 -11748 -15880
rect -12548 -16640 -11748 -16600
rect -11136 -15880 -10336 -15840
rect -11136 -16600 -11096 -15880
rect -10376 -16600 -10336 -15880
rect -11136 -16640 -10336 -16600
rect -9724 -15880 -8924 -15840
rect -9724 -16600 -9684 -15880
rect -8964 -16600 -8924 -15880
rect -9724 -16640 -8924 -16600
rect -8312 -15880 -7512 -15840
rect -8312 -16600 -8272 -15880
rect -7552 -16600 -7512 -15880
rect -8312 -16640 -7512 -16600
rect -6900 -15880 -6100 -15840
rect -6900 -16600 -6860 -15880
rect -6140 -16600 -6100 -15880
rect -6900 -16640 -6100 -16600
rect -5488 -15880 -4688 -15840
rect -5488 -16600 -5448 -15880
rect -4728 -16600 -4688 -15880
rect -5488 -16640 -4688 -16600
rect -4076 -15880 -3276 -15840
rect -4076 -16600 -4036 -15880
rect -3316 -16600 -3276 -15880
rect -4076 -16640 -3276 -16600
rect -2664 -15880 -1864 -15840
rect -2664 -16600 -2624 -15880
rect -1904 -16600 -1864 -15880
rect -2664 -16640 -1864 -16600
rect -1252 -15880 -452 -15840
rect -1252 -16600 -1212 -15880
rect -492 -16600 -452 -15880
rect -1252 -16640 -452 -16600
rect 160 -15880 960 -15840
rect 160 -16600 200 -15880
rect 920 -16600 960 -15880
rect 160 -16640 960 -16600
rect 1572 -15880 2372 -15840
rect 1572 -16600 1612 -15880
rect 2332 -16600 2372 -15880
rect 1572 -16640 2372 -16600
rect 2984 -15880 3784 -15840
rect 2984 -16600 3024 -15880
rect 3744 -16600 3784 -15880
rect 2984 -16640 3784 -16600
rect 4396 -15880 5196 -15840
rect 4396 -16600 4436 -15880
rect 5156 -16600 5196 -15880
rect 4396 -16640 5196 -16600
rect 5808 -15880 6608 -15840
rect 5808 -16600 5848 -15880
rect 6568 -16600 6608 -15880
rect 5808 -16640 6608 -16600
rect 7220 -15880 8020 -15840
rect 7220 -16600 7260 -15880
rect 7980 -16600 8020 -15880
rect 7220 -16640 8020 -16600
rect 8632 -15880 9432 -15840
rect 8632 -16600 8672 -15880
rect 9392 -16600 9432 -15880
rect 8632 -16640 9432 -16600
rect 10044 -15880 10844 -15840
rect 10044 -16600 10084 -15880
rect 10804 -16600 10844 -15880
rect 10044 -16640 10844 -16600
rect 11456 -15880 12256 -15840
rect 11456 -16600 11496 -15880
rect 12216 -16600 12256 -15880
rect 11456 -16640 12256 -16600
rect 12868 -15880 13668 -15840
rect 12868 -16600 12908 -15880
rect 13628 -16600 13668 -15880
rect 12868 -16640 13668 -16600
rect 14280 -15880 15080 -15840
rect 14280 -16600 14320 -15880
rect 15040 -16600 15080 -15880
rect 14280 -16640 15080 -16600
rect 15692 -15880 16492 -15840
rect 15692 -16600 15732 -15880
rect 16452 -16600 16492 -15880
rect 15692 -16640 16492 -16600
rect 17104 -15880 17904 -15840
rect 17104 -16600 17144 -15880
rect 17864 -16600 17904 -15880
rect 17104 -16640 17904 -16600
rect 18516 -15880 19316 -15840
rect 18516 -16600 18556 -15880
rect 19276 -16600 19316 -15880
rect 18516 -16640 19316 -16600
rect 19928 -15880 20728 -15840
rect 19928 -16600 19968 -15880
rect 20688 -16600 20728 -15880
rect 19928 -16640 20728 -16600
rect 21340 -15880 22140 -15840
rect 21340 -16600 21380 -15880
rect 22100 -16600 22140 -15880
rect 21340 -16640 22140 -16600
rect 22752 -15880 23552 -15840
rect 22752 -16600 22792 -15880
rect 23512 -16600 23552 -15880
rect 22752 -16640 23552 -16600
rect -23844 -17000 -23044 -16960
rect -23844 -17720 -23804 -17000
rect -23084 -17720 -23044 -17000
rect -23844 -17760 -23044 -17720
rect -22432 -17000 -21632 -16960
rect -22432 -17720 -22392 -17000
rect -21672 -17720 -21632 -17000
rect -22432 -17760 -21632 -17720
rect -21020 -17000 -20220 -16960
rect -21020 -17720 -20980 -17000
rect -20260 -17720 -20220 -17000
rect -21020 -17760 -20220 -17720
rect -19608 -17000 -18808 -16960
rect -19608 -17720 -19568 -17000
rect -18848 -17720 -18808 -17000
rect -19608 -17760 -18808 -17720
rect -18196 -17000 -17396 -16960
rect -18196 -17720 -18156 -17000
rect -17436 -17720 -17396 -17000
rect -18196 -17760 -17396 -17720
rect -16784 -17000 -15984 -16960
rect -16784 -17720 -16744 -17000
rect -16024 -17720 -15984 -17000
rect -16784 -17760 -15984 -17720
rect -15372 -17000 -14572 -16960
rect -15372 -17720 -15332 -17000
rect -14612 -17720 -14572 -17000
rect -15372 -17760 -14572 -17720
rect -13960 -17000 -13160 -16960
rect -13960 -17720 -13920 -17000
rect -13200 -17720 -13160 -17000
rect -13960 -17760 -13160 -17720
rect -12548 -17000 -11748 -16960
rect -12548 -17720 -12508 -17000
rect -11788 -17720 -11748 -17000
rect -12548 -17760 -11748 -17720
rect -11136 -17000 -10336 -16960
rect -11136 -17720 -11096 -17000
rect -10376 -17720 -10336 -17000
rect -11136 -17760 -10336 -17720
rect -9724 -17000 -8924 -16960
rect -9724 -17720 -9684 -17000
rect -8964 -17720 -8924 -17000
rect -9724 -17760 -8924 -17720
rect -8312 -17000 -7512 -16960
rect -8312 -17720 -8272 -17000
rect -7552 -17720 -7512 -17000
rect -8312 -17760 -7512 -17720
rect -6900 -17000 -6100 -16960
rect -6900 -17720 -6860 -17000
rect -6140 -17720 -6100 -17000
rect -6900 -17760 -6100 -17720
rect -5488 -17000 -4688 -16960
rect -5488 -17720 -5448 -17000
rect -4728 -17720 -4688 -17000
rect -5488 -17760 -4688 -17720
rect -4076 -17000 -3276 -16960
rect -4076 -17720 -4036 -17000
rect -3316 -17720 -3276 -17000
rect -4076 -17760 -3276 -17720
rect -2664 -17000 -1864 -16960
rect -2664 -17720 -2624 -17000
rect -1904 -17720 -1864 -17000
rect -2664 -17760 -1864 -17720
rect -1252 -17000 -452 -16960
rect -1252 -17720 -1212 -17000
rect -492 -17720 -452 -17000
rect -1252 -17760 -452 -17720
rect 160 -17000 960 -16960
rect 160 -17720 200 -17000
rect 920 -17720 960 -17000
rect 160 -17760 960 -17720
rect 1572 -17000 2372 -16960
rect 1572 -17720 1612 -17000
rect 2332 -17720 2372 -17000
rect 1572 -17760 2372 -17720
rect 2984 -17000 3784 -16960
rect 2984 -17720 3024 -17000
rect 3744 -17720 3784 -17000
rect 2984 -17760 3784 -17720
rect 4396 -17000 5196 -16960
rect 4396 -17720 4436 -17000
rect 5156 -17720 5196 -17000
rect 4396 -17760 5196 -17720
rect 5808 -17000 6608 -16960
rect 5808 -17720 5848 -17000
rect 6568 -17720 6608 -17000
rect 5808 -17760 6608 -17720
rect 7220 -17000 8020 -16960
rect 7220 -17720 7260 -17000
rect 7980 -17720 8020 -17000
rect 7220 -17760 8020 -17720
rect 8632 -17000 9432 -16960
rect 8632 -17720 8672 -17000
rect 9392 -17720 9432 -17000
rect 8632 -17760 9432 -17720
rect 10044 -17000 10844 -16960
rect 10044 -17720 10084 -17000
rect 10804 -17720 10844 -17000
rect 10044 -17760 10844 -17720
rect 11456 -17000 12256 -16960
rect 11456 -17720 11496 -17000
rect 12216 -17720 12256 -17000
rect 11456 -17760 12256 -17720
rect 12868 -17000 13668 -16960
rect 12868 -17720 12908 -17000
rect 13628 -17720 13668 -17000
rect 12868 -17760 13668 -17720
rect 14280 -17000 15080 -16960
rect 14280 -17720 14320 -17000
rect 15040 -17720 15080 -17000
rect 14280 -17760 15080 -17720
rect 15692 -17000 16492 -16960
rect 15692 -17720 15732 -17000
rect 16452 -17720 16492 -17000
rect 15692 -17760 16492 -17720
rect 17104 -17000 17904 -16960
rect 17104 -17720 17144 -17000
rect 17864 -17720 17904 -17000
rect 17104 -17760 17904 -17720
rect 18516 -17000 19316 -16960
rect 18516 -17720 18556 -17000
rect 19276 -17720 19316 -17000
rect 18516 -17760 19316 -17720
rect 19928 -17000 20728 -16960
rect 19928 -17720 19968 -17000
rect 20688 -17720 20728 -17000
rect 19928 -17760 20728 -17720
rect 21340 -17000 22140 -16960
rect 21340 -17720 21380 -17000
rect 22100 -17720 22140 -17000
rect 21340 -17760 22140 -17720
rect 22752 -17000 23552 -16960
rect 22752 -17720 22792 -17000
rect 23512 -17720 23552 -17000
rect 22752 -17760 23552 -17720
rect -23844 -18120 -23044 -18080
rect -23844 -18840 -23804 -18120
rect -23084 -18840 -23044 -18120
rect -23844 -18880 -23044 -18840
rect -22432 -18120 -21632 -18080
rect -22432 -18840 -22392 -18120
rect -21672 -18840 -21632 -18120
rect -22432 -18880 -21632 -18840
rect -21020 -18120 -20220 -18080
rect -21020 -18840 -20980 -18120
rect -20260 -18840 -20220 -18120
rect -21020 -18880 -20220 -18840
rect -19608 -18120 -18808 -18080
rect -19608 -18840 -19568 -18120
rect -18848 -18840 -18808 -18120
rect -19608 -18880 -18808 -18840
rect -18196 -18120 -17396 -18080
rect -18196 -18840 -18156 -18120
rect -17436 -18840 -17396 -18120
rect -18196 -18880 -17396 -18840
rect -16784 -18120 -15984 -18080
rect -16784 -18840 -16744 -18120
rect -16024 -18840 -15984 -18120
rect -16784 -18880 -15984 -18840
rect -15372 -18120 -14572 -18080
rect -15372 -18840 -15332 -18120
rect -14612 -18840 -14572 -18120
rect -15372 -18880 -14572 -18840
rect -13960 -18120 -13160 -18080
rect -13960 -18840 -13920 -18120
rect -13200 -18840 -13160 -18120
rect -13960 -18880 -13160 -18840
rect -12548 -18120 -11748 -18080
rect -12548 -18840 -12508 -18120
rect -11788 -18840 -11748 -18120
rect -12548 -18880 -11748 -18840
rect -11136 -18120 -10336 -18080
rect -11136 -18840 -11096 -18120
rect -10376 -18840 -10336 -18120
rect -11136 -18880 -10336 -18840
rect -9724 -18120 -8924 -18080
rect -9724 -18840 -9684 -18120
rect -8964 -18840 -8924 -18120
rect -9724 -18880 -8924 -18840
rect -8312 -18120 -7512 -18080
rect -8312 -18840 -8272 -18120
rect -7552 -18840 -7512 -18120
rect -8312 -18880 -7512 -18840
rect -6900 -18120 -6100 -18080
rect -6900 -18840 -6860 -18120
rect -6140 -18840 -6100 -18120
rect -6900 -18880 -6100 -18840
rect -5488 -18120 -4688 -18080
rect -5488 -18840 -5448 -18120
rect -4728 -18840 -4688 -18120
rect -5488 -18880 -4688 -18840
rect -4076 -18120 -3276 -18080
rect -4076 -18840 -4036 -18120
rect -3316 -18840 -3276 -18120
rect -4076 -18880 -3276 -18840
rect -2664 -18120 -1864 -18080
rect -2664 -18840 -2624 -18120
rect -1904 -18840 -1864 -18120
rect -2664 -18880 -1864 -18840
rect -1252 -18120 -452 -18080
rect -1252 -18840 -1212 -18120
rect -492 -18840 -452 -18120
rect -1252 -18880 -452 -18840
rect 160 -18120 960 -18080
rect 160 -18840 200 -18120
rect 920 -18840 960 -18120
rect 160 -18880 960 -18840
rect 1572 -18120 2372 -18080
rect 1572 -18840 1612 -18120
rect 2332 -18840 2372 -18120
rect 1572 -18880 2372 -18840
rect 2984 -18120 3784 -18080
rect 2984 -18840 3024 -18120
rect 3744 -18840 3784 -18120
rect 2984 -18880 3784 -18840
rect 4396 -18120 5196 -18080
rect 4396 -18840 4436 -18120
rect 5156 -18840 5196 -18120
rect 4396 -18880 5196 -18840
rect 5808 -18120 6608 -18080
rect 5808 -18840 5848 -18120
rect 6568 -18840 6608 -18120
rect 5808 -18880 6608 -18840
rect 7220 -18120 8020 -18080
rect 7220 -18840 7260 -18120
rect 7980 -18840 8020 -18120
rect 7220 -18880 8020 -18840
rect 8632 -18120 9432 -18080
rect 8632 -18840 8672 -18120
rect 9392 -18840 9432 -18120
rect 8632 -18880 9432 -18840
rect 10044 -18120 10844 -18080
rect 10044 -18840 10084 -18120
rect 10804 -18840 10844 -18120
rect 10044 -18880 10844 -18840
rect 11456 -18120 12256 -18080
rect 11456 -18840 11496 -18120
rect 12216 -18840 12256 -18120
rect 11456 -18880 12256 -18840
rect 12868 -18120 13668 -18080
rect 12868 -18840 12908 -18120
rect 13628 -18840 13668 -18120
rect 12868 -18880 13668 -18840
rect 14280 -18120 15080 -18080
rect 14280 -18840 14320 -18120
rect 15040 -18840 15080 -18120
rect 14280 -18880 15080 -18840
rect 15692 -18120 16492 -18080
rect 15692 -18840 15732 -18120
rect 16452 -18840 16492 -18120
rect 15692 -18880 16492 -18840
rect 17104 -18120 17904 -18080
rect 17104 -18840 17144 -18120
rect 17864 -18840 17904 -18120
rect 17104 -18880 17904 -18840
rect 18516 -18120 19316 -18080
rect 18516 -18840 18556 -18120
rect 19276 -18840 19316 -18120
rect 18516 -18880 19316 -18840
rect 19928 -18120 20728 -18080
rect 19928 -18840 19968 -18120
rect 20688 -18840 20728 -18120
rect 19928 -18880 20728 -18840
rect 21340 -18120 22140 -18080
rect 21340 -18840 21380 -18120
rect 22100 -18840 22140 -18120
rect 21340 -18880 22140 -18840
rect 22752 -18120 23552 -18080
rect 22752 -18840 22792 -18120
rect 23512 -18840 23552 -18120
rect 22752 -18880 23552 -18840
<< mimcapcontact >>
rect -23804 18120 -23084 18840
rect -22392 18120 -21672 18840
rect -20980 18120 -20260 18840
rect -19568 18120 -18848 18840
rect -18156 18120 -17436 18840
rect -16744 18120 -16024 18840
rect -15332 18120 -14612 18840
rect -13920 18120 -13200 18840
rect -12508 18120 -11788 18840
rect -11096 18120 -10376 18840
rect -9684 18120 -8964 18840
rect -8272 18120 -7552 18840
rect -6860 18120 -6140 18840
rect -5448 18120 -4728 18840
rect -4036 18120 -3316 18840
rect -2624 18120 -1904 18840
rect -1212 18120 -492 18840
rect 200 18120 920 18840
rect 1612 18120 2332 18840
rect 3024 18120 3744 18840
rect 4436 18120 5156 18840
rect 5848 18120 6568 18840
rect 7260 18120 7980 18840
rect 8672 18120 9392 18840
rect 10084 18120 10804 18840
rect 11496 18120 12216 18840
rect 12908 18120 13628 18840
rect 14320 18120 15040 18840
rect 15732 18120 16452 18840
rect 17144 18120 17864 18840
rect 18556 18120 19276 18840
rect 19968 18120 20688 18840
rect 21380 18120 22100 18840
rect 22792 18120 23512 18840
rect -23804 17000 -23084 17720
rect -22392 17000 -21672 17720
rect -20980 17000 -20260 17720
rect -19568 17000 -18848 17720
rect -18156 17000 -17436 17720
rect -16744 17000 -16024 17720
rect -15332 17000 -14612 17720
rect -13920 17000 -13200 17720
rect -12508 17000 -11788 17720
rect -11096 17000 -10376 17720
rect -9684 17000 -8964 17720
rect -8272 17000 -7552 17720
rect -6860 17000 -6140 17720
rect -5448 17000 -4728 17720
rect -4036 17000 -3316 17720
rect -2624 17000 -1904 17720
rect -1212 17000 -492 17720
rect 200 17000 920 17720
rect 1612 17000 2332 17720
rect 3024 17000 3744 17720
rect 4436 17000 5156 17720
rect 5848 17000 6568 17720
rect 7260 17000 7980 17720
rect 8672 17000 9392 17720
rect 10084 17000 10804 17720
rect 11496 17000 12216 17720
rect 12908 17000 13628 17720
rect 14320 17000 15040 17720
rect 15732 17000 16452 17720
rect 17144 17000 17864 17720
rect 18556 17000 19276 17720
rect 19968 17000 20688 17720
rect 21380 17000 22100 17720
rect 22792 17000 23512 17720
rect -23804 15880 -23084 16600
rect -22392 15880 -21672 16600
rect -20980 15880 -20260 16600
rect -19568 15880 -18848 16600
rect -18156 15880 -17436 16600
rect -16744 15880 -16024 16600
rect -15332 15880 -14612 16600
rect -13920 15880 -13200 16600
rect -12508 15880 -11788 16600
rect -11096 15880 -10376 16600
rect -9684 15880 -8964 16600
rect -8272 15880 -7552 16600
rect -6860 15880 -6140 16600
rect -5448 15880 -4728 16600
rect -4036 15880 -3316 16600
rect -2624 15880 -1904 16600
rect -1212 15880 -492 16600
rect 200 15880 920 16600
rect 1612 15880 2332 16600
rect 3024 15880 3744 16600
rect 4436 15880 5156 16600
rect 5848 15880 6568 16600
rect 7260 15880 7980 16600
rect 8672 15880 9392 16600
rect 10084 15880 10804 16600
rect 11496 15880 12216 16600
rect 12908 15880 13628 16600
rect 14320 15880 15040 16600
rect 15732 15880 16452 16600
rect 17144 15880 17864 16600
rect 18556 15880 19276 16600
rect 19968 15880 20688 16600
rect 21380 15880 22100 16600
rect 22792 15880 23512 16600
rect -23804 14760 -23084 15480
rect -22392 14760 -21672 15480
rect -20980 14760 -20260 15480
rect -19568 14760 -18848 15480
rect -18156 14760 -17436 15480
rect -16744 14760 -16024 15480
rect -15332 14760 -14612 15480
rect -13920 14760 -13200 15480
rect -12508 14760 -11788 15480
rect -11096 14760 -10376 15480
rect -9684 14760 -8964 15480
rect -8272 14760 -7552 15480
rect -6860 14760 -6140 15480
rect -5448 14760 -4728 15480
rect -4036 14760 -3316 15480
rect -2624 14760 -1904 15480
rect -1212 14760 -492 15480
rect 200 14760 920 15480
rect 1612 14760 2332 15480
rect 3024 14760 3744 15480
rect 4436 14760 5156 15480
rect 5848 14760 6568 15480
rect 7260 14760 7980 15480
rect 8672 14760 9392 15480
rect 10084 14760 10804 15480
rect 11496 14760 12216 15480
rect 12908 14760 13628 15480
rect 14320 14760 15040 15480
rect 15732 14760 16452 15480
rect 17144 14760 17864 15480
rect 18556 14760 19276 15480
rect 19968 14760 20688 15480
rect 21380 14760 22100 15480
rect 22792 14760 23512 15480
rect -23804 13640 -23084 14360
rect -22392 13640 -21672 14360
rect -20980 13640 -20260 14360
rect -19568 13640 -18848 14360
rect -18156 13640 -17436 14360
rect -16744 13640 -16024 14360
rect -15332 13640 -14612 14360
rect -13920 13640 -13200 14360
rect -12508 13640 -11788 14360
rect -11096 13640 -10376 14360
rect -9684 13640 -8964 14360
rect -8272 13640 -7552 14360
rect -6860 13640 -6140 14360
rect -5448 13640 -4728 14360
rect -4036 13640 -3316 14360
rect -2624 13640 -1904 14360
rect -1212 13640 -492 14360
rect 200 13640 920 14360
rect 1612 13640 2332 14360
rect 3024 13640 3744 14360
rect 4436 13640 5156 14360
rect 5848 13640 6568 14360
rect 7260 13640 7980 14360
rect 8672 13640 9392 14360
rect 10084 13640 10804 14360
rect 11496 13640 12216 14360
rect 12908 13640 13628 14360
rect 14320 13640 15040 14360
rect 15732 13640 16452 14360
rect 17144 13640 17864 14360
rect 18556 13640 19276 14360
rect 19968 13640 20688 14360
rect 21380 13640 22100 14360
rect 22792 13640 23512 14360
rect -23804 12520 -23084 13240
rect -22392 12520 -21672 13240
rect -20980 12520 -20260 13240
rect -19568 12520 -18848 13240
rect -18156 12520 -17436 13240
rect -16744 12520 -16024 13240
rect -15332 12520 -14612 13240
rect -13920 12520 -13200 13240
rect -12508 12520 -11788 13240
rect -11096 12520 -10376 13240
rect -9684 12520 -8964 13240
rect -8272 12520 -7552 13240
rect -6860 12520 -6140 13240
rect -5448 12520 -4728 13240
rect -4036 12520 -3316 13240
rect -2624 12520 -1904 13240
rect -1212 12520 -492 13240
rect 200 12520 920 13240
rect 1612 12520 2332 13240
rect 3024 12520 3744 13240
rect 4436 12520 5156 13240
rect 5848 12520 6568 13240
rect 7260 12520 7980 13240
rect 8672 12520 9392 13240
rect 10084 12520 10804 13240
rect 11496 12520 12216 13240
rect 12908 12520 13628 13240
rect 14320 12520 15040 13240
rect 15732 12520 16452 13240
rect 17144 12520 17864 13240
rect 18556 12520 19276 13240
rect 19968 12520 20688 13240
rect 21380 12520 22100 13240
rect 22792 12520 23512 13240
rect -23804 11400 -23084 12120
rect -22392 11400 -21672 12120
rect -20980 11400 -20260 12120
rect -19568 11400 -18848 12120
rect -18156 11400 -17436 12120
rect -16744 11400 -16024 12120
rect -15332 11400 -14612 12120
rect -13920 11400 -13200 12120
rect -12508 11400 -11788 12120
rect -11096 11400 -10376 12120
rect -9684 11400 -8964 12120
rect -8272 11400 -7552 12120
rect -6860 11400 -6140 12120
rect -5448 11400 -4728 12120
rect -4036 11400 -3316 12120
rect -2624 11400 -1904 12120
rect -1212 11400 -492 12120
rect 200 11400 920 12120
rect 1612 11400 2332 12120
rect 3024 11400 3744 12120
rect 4436 11400 5156 12120
rect 5848 11400 6568 12120
rect 7260 11400 7980 12120
rect 8672 11400 9392 12120
rect 10084 11400 10804 12120
rect 11496 11400 12216 12120
rect 12908 11400 13628 12120
rect 14320 11400 15040 12120
rect 15732 11400 16452 12120
rect 17144 11400 17864 12120
rect 18556 11400 19276 12120
rect 19968 11400 20688 12120
rect 21380 11400 22100 12120
rect 22792 11400 23512 12120
rect -23804 10280 -23084 11000
rect -22392 10280 -21672 11000
rect -20980 10280 -20260 11000
rect -19568 10280 -18848 11000
rect -18156 10280 -17436 11000
rect -16744 10280 -16024 11000
rect -15332 10280 -14612 11000
rect -13920 10280 -13200 11000
rect -12508 10280 -11788 11000
rect -11096 10280 -10376 11000
rect -9684 10280 -8964 11000
rect -8272 10280 -7552 11000
rect -6860 10280 -6140 11000
rect -5448 10280 -4728 11000
rect -4036 10280 -3316 11000
rect -2624 10280 -1904 11000
rect -1212 10280 -492 11000
rect 200 10280 920 11000
rect 1612 10280 2332 11000
rect 3024 10280 3744 11000
rect 4436 10280 5156 11000
rect 5848 10280 6568 11000
rect 7260 10280 7980 11000
rect 8672 10280 9392 11000
rect 10084 10280 10804 11000
rect 11496 10280 12216 11000
rect 12908 10280 13628 11000
rect 14320 10280 15040 11000
rect 15732 10280 16452 11000
rect 17144 10280 17864 11000
rect 18556 10280 19276 11000
rect 19968 10280 20688 11000
rect 21380 10280 22100 11000
rect 22792 10280 23512 11000
rect -23804 9160 -23084 9880
rect -22392 9160 -21672 9880
rect -20980 9160 -20260 9880
rect -19568 9160 -18848 9880
rect -18156 9160 -17436 9880
rect -16744 9160 -16024 9880
rect -15332 9160 -14612 9880
rect -13920 9160 -13200 9880
rect -12508 9160 -11788 9880
rect -11096 9160 -10376 9880
rect -9684 9160 -8964 9880
rect -8272 9160 -7552 9880
rect -6860 9160 -6140 9880
rect -5448 9160 -4728 9880
rect -4036 9160 -3316 9880
rect -2624 9160 -1904 9880
rect -1212 9160 -492 9880
rect 200 9160 920 9880
rect 1612 9160 2332 9880
rect 3024 9160 3744 9880
rect 4436 9160 5156 9880
rect 5848 9160 6568 9880
rect 7260 9160 7980 9880
rect 8672 9160 9392 9880
rect 10084 9160 10804 9880
rect 11496 9160 12216 9880
rect 12908 9160 13628 9880
rect 14320 9160 15040 9880
rect 15732 9160 16452 9880
rect 17144 9160 17864 9880
rect 18556 9160 19276 9880
rect 19968 9160 20688 9880
rect 21380 9160 22100 9880
rect 22792 9160 23512 9880
rect -23804 8040 -23084 8760
rect -22392 8040 -21672 8760
rect -20980 8040 -20260 8760
rect -19568 8040 -18848 8760
rect -18156 8040 -17436 8760
rect -16744 8040 -16024 8760
rect -15332 8040 -14612 8760
rect -13920 8040 -13200 8760
rect -12508 8040 -11788 8760
rect -11096 8040 -10376 8760
rect -9684 8040 -8964 8760
rect -8272 8040 -7552 8760
rect -6860 8040 -6140 8760
rect -5448 8040 -4728 8760
rect -4036 8040 -3316 8760
rect -2624 8040 -1904 8760
rect -1212 8040 -492 8760
rect 200 8040 920 8760
rect 1612 8040 2332 8760
rect 3024 8040 3744 8760
rect 4436 8040 5156 8760
rect 5848 8040 6568 8760
rect 7260 8040 7980 8760
rect 8672 8040 9392 8760
rect 10084 8040 10804 8760
rect 11496 8040 12216 8760
rect 12908 8040 13628 8760
rect 14320 8040 15040 8760
rect 15732 8040 16452 8760
rect 17144 8040 17864 8760
rect 18556 8040 19276 8760
rect 19968 8040 20688 8760
rect 21380 8040 22100 8760
rect 22792 8040 23512 8760
rect -23804 6920 -23084 7640
rect -22392 6920 -21672 7640
rect -20980 6920 -20260 7640
rect -19568 6920 -18848 7640
rect -18156 6920 -17436 7640
rect -16744 6920 -16024 7640
rect -15332 6920 -14612 7640
rect -13920 6920 -13200 7640
rect -12508 6920 -11788 7640
rect -11096 6920 -10376 7640
rect -9684 6920 -8964 7640
rect -8272 6920 -7552 7640
rect -6860 6920 -6140 7640
rect -5448 6920 -4728 7640
rect -4036 6920 -3316 7640
rect -2624 6920 -1904 7640
rect -1212 6920 -492 7640
rect 200 6920 920 7640
rect 1612 6920 2332 7640
rect 3024 6920 3744 7640
rect 4436 6920 5156 7640
rect 5848 6920 6568 7640
rect 7260 6920 7980 7640
rect 8672 6920 9392 7640
rect 10084 6920 10804 7640
rect 11496 6920 12216 7640
rect 12908 6920 13628 7640
rect 14320 6920 15040 7640
rect 15732 6920 16452 7640
rect 17144 6920 17864 7640
rect 18556 6920 19276 7640
rect 19968 6920 20688 7640
rect 21380 6920 22100 7640
rect 22792 6920 23512 7640
rect -23804 5800 -23084 6520
rect -22392 5800 -21672 6520
rect -20980 5800 -20260 6520
rect -19568 5800 -18848 6520
rect -18156 5800 -17436 6520
rect -16744 5800 -16024 6520
rect -15332 5800 -14612 6520
rect -13920 5800 -13200 6520
rect -12508 5800 -11788 6520
rect -11096 5800 -10376 6520
rect -9684 5800 -8964 6520
rect -8272 5800 -7552 6520
rect -6860 5800 -6140 6520
rect -5448 5800 -4728 6520
rect -4036 5800 -3316 6520
rect -2624 5800 -1904 6520
rect -1212 5800 -492 6520
rect 200 5800 920 6520
rect 1612 5800 2332 6520
rect 3024 5800 3744 6520
rect 4436 5800 5156 6520
rect 5848 5800 6568 6520
rect 7260 5800 7980 6520
rect 8672 5800 9392 6520
rect 10084 5800 10804 6520
rect 11496 5800 12216 6520
rect 12908 5800 13628 6520
rect 14320 5800 15040 6520
rect 15732 5800 16452 6520
rect 17144 5800 17864 6520
rect 18556 5800 19276 6520
rect 19968 5800 20688 6520
rect 21380 5800 22100 6520
rect 22792 5800 23512 6520
rect -23804 4680 -23084 5400
rect -22392 4680 -21672 5400
rect -20980 4680 -20260 5400
rect -19568 4680 -18848 5400
rect -18156 4680 -17436 5400
rect -16744 4680 -16024 5400
rect -15332 4680 -14612 5400
rect -13920 4680 -13200 5400
rect -12508 4680 -11788 5400
rect -11096 4680 -10376 5400
rect -9684 4680 -8964 5400
rect -8272 4680 -7552 5400
rect -6860 4680 -6140 5400
rect -5448 4680 -4728 5400
rect -4036 4680 -3316 5400
rect -2624 4680 -1904 5400
rect -1212 4680 -492 5400
rect 200 4680 920 5400
rect 1612 4680 2332 5400
rect 3024 4680 3744 5400
rect 4436 4680 5156 5400
rect 5848 4680 6568 5400
rect 7260 4680 7980 5400
rect 8672 4680 9392 5400
rect 10084 4680 10804 5400
rect 11496 4680 12216 5400
rect 12908 4680 13628 5400
rect 14320 4680 15040 5400
rect 15732 4680 16452 5400
rect 17144 4680 17864 5400
rect 18556 4680 19276 5400
rect 19968 4680 20688 5400
rect 21380 4680 22100 5400
rect 22792 4680 23512 5400
rect -23804 3560 -23084 4280
rect -22392 3560 -21672 4280
rect -20980 3560 -20260 4280
rect -19568 3560 -18848 4280
rect -18156 3560 -17436 4280
rect -16744 3560 -16024 4280
rect -15332 3560 -14612 4280
rect -13920 3560 -13200 4280
rect -12508 3560 -11788 4280
rect -11096 3560 -10376 4280
rect -9684 3560 -8964 4280
rect -8272 3560 -7552 4280
rect -6860 3560 -6140 4280
rect -5448 3560 -4728 4280
rect -4036 3560 -3316 4280
rect -2624 3560 -1904 4280
rect -1212 3560 -492 4280
rect 200 3560 920 4280
rect 1612 3560 2332 4280
rect 3024 3560 3744 4280
rect 4436 3560 5156 4280
rect 5848 3560 6568 4280
rect 7260 3560 7980 4280
rect 8672 3560 9392 4280
rect 10084 3560 10804 4280
rect 11496 3560 12216 4280
rect 12908 3560 13628 4280
rect 14320 3560 15040 4280
rect 15732 3560 16452 4280
rect 17144 3560 17864 4280
rect 18556 3560 19276 4280
rect 19968 3560 20688 4280
rect 21380 3560 22100 4280
rect 22792 3560 23512 4280
rect -23804 2440 -23084 3160
rect -22392 2440 -21672 3160
rect -20980 2440 -20260 3160
rect -19568 2440 -18848 3160
rect -18156 2440 -17436 3160
rect -16744 2440 -16024 3160
rect -15332 2440 -14612 3160
rect -13920 2440 -13200 3160
rect -12508 2440 -11788 3160
rect -11096 2440 -10376 3160
rect -9684 2440 -8964 3160
rect -8272 2440 -7552 3160
rect -6860 2440 -6140 3160
rect -5448 2440 -4728 3160
rect -4036 2440 -3316 3160
rect -2624 2440 -1904 3160
rect -1212 2440 -492 3160
rect 200 2440 920 3160
rect 1612 2440 2332 3160
rect 3024 2440 3744 3160
rect 4436 2440 5156 3160
rect 5848 2440 6568 3160
rect 7260 2440 7980 3160
rect 8672 2440 9392 3160
rect 10084 2440 10804 3160
rect 11496 2440 12216 3160
rect 12908 2440 13628 3160
rect 14320 2440 15040 3160
rect 15732 2440 16452 3160
rect 17144 2440 17864 3160
rect 18556 2440 19276 3160
rect 19968 2440 20688 3160
rect 21380 2440 22100 3160
rect 22792 2440 23512 3160
rect -23804 1320 -23084 2040
rect -22392 1320 -21672 2040
rect -20980 1320 -20260 2040
rect -19568 1320 -18848 2040
rect -18156 1320 -17436 2040
rect -16744 1320 -16024 2040
rect -15332 1320 -14612 2040
rect -13920 1320 -13200 2040
rect -12508 1320 -11788 2040
rect -11096 1320 -10376 2040
rect -9684 1320 -8964 2040
rect -8272 1320 -7552 2040
rect -6860 1320 -6140 2040
rect -5448 1320 -4728 2040
rect -4036 1320 -3316 2040
rect -2624 1320 -1904 2040
rect -1212 1320 -492 2040
rect 200 1320 920 2040
rect 1612 1320 2332 2040
rect 3024 1320 3744 2040
rect 4436 1320 5156 2040
rect 5848 1320 6568 2040
rect 7260 1320 7980 2040
rect 8672 1320 9392 2040
rect 10084 1320 10804 2040
rect 11496 1320 12216 2040
rect 12908 1320 13628 2040
rect 14320 1320 15040 2040
rect 15732 1320 16452 2040
rect 17144 1320 17864 2040
rect 18556 1320 19276 2040
rect 19968 1320 20688 2040
rect 21380 1320 22100 2040
rect 22792 1320 23512 2040
rect -23804 200 -23084 920
rect -22392 200 -21672 920
rect -20980 200 -20260 920
rect -19568 200 -18848 920
rect -18156 200 -17436 920
rect -16744 200 -16024 920
rect -15332 200 -14612 920
rect -13920 200 -13200 920
rect -12508 200 -11788 920
rect -11096 200 -10376 920
rect -9684 200 -8964 920
rect -8272 200 -7552 920
rect -6860 200 -6140 920
rect -5448 200 -4728 920
rect -4036 200 -3316 920
rect -2624 200 -1904 920
rect -1212 200 -492 920
rect 200 200 920 920
rect 1612 200 2332 920
rect 3024 200 3744 920
rect 4436 200 5156 920
rect 5848 200 6568 920
rect 7260 200 7980 920
rect 8672 200 9392 920
rect 10084 200 10804 920
rect 11496 200 12216 920
rect 12908 200 13628 920
rect 14320 200 15040 920
rect 15732 200 16452 920
rect 17144 200 17864 920
rect 18556 200 19276 920
rect 19968 200 20688 920
rect 21380 200 22100 920
rect 22792 200 23512 920
rect -23804 -920 -23084 -200
rect -22392 -920 -21672 -200
rect -20980 -920 -20260 -200
rect -19568 -920 -18848 -200
rect -18156 -920 -17436 -200
rect -16744 -920 -16024 -200
rect -15332 -920 -14612 -200
rect -13920 -920 -13200 -200
rect -12508 -920 -11788 -200
rect -11096 -920 -10376 -200
rect -9684 -920 -8964 -200
rect -8272 -920 -7552 -200
rect -6860 -920 -6140 -200
rect -5448 -920 -4728 -200
rect -4036 -920 -3316 -200
rect -2624 -920 -1904 -200
rect -1212 -920 -492 -200
rect 200 -920 920 -200
rect 1612 -920 2332 -200
rect 3024 -920 3744 -200
rect 4436 -920 5156 -200
rect 5848 -920 6568 -200
rect 7260 -920 7980 -200
rect 8672 -920 9392 -200
rect 10084 -920 10804 -200
rect 11496 -920 12216 -200
rect 12908 -920 13628 -200
rect 14320 -920 15040 -200
rect 15732 -920 16452 -200
rect 17144 -920 17864 -200
rect 18556 -920 19276 -200
rect 19968 -920 20688 -200
rect 21380 -920 22100 -200
rect 22792 -920 23512 -200
rect -23804 -2040 -23084 -1320
rect -22392 -2040 -21672 -1320
rect -20980 -2040 -20260 -1320
rect -19568 -2040 -18848 -1320
rect -18156 -2040 -17436 -1320
rect -16744 -2040 -16024 -1320
rect -15332 -2040 -14612 -1320
rect -13920 -2040 -13200 -1320
rect -12508 -2040 -11788 -1320
rect -11096 -2040 -10376 -1320
rect -9684 -2040 -8964 -1320
rect -8272 -2040 -7552 -1320
rect -6860 -2040 -6140 -1320
rect -5448 -2040 -4728 -1320
rect -4036 -2040 -3316 -1320
rect -2624 -2040 -1904 -1320
rect -1212 -2040 -492 -1320
rect 200 -2040 920 -1320
rect 1612 -2040 2332 -1320
rect 3024 -2040 3744 -1320
rect 4436 -2040 5156 -1320
rect 5848 -2040 6568 -1320
rect 7260 -2040 7980 -1320
rect 8672 -2040 9392 -1320
rect 10084 -2040 10804 -1320
rect 11496 -2040 12216 -1320
rect 12908 -2040 13628 -1320
rect 14320 -2040 15040 -1320
rect 15732 -2040 16452 -1320
rect 17144 -2040 17864 -1320
rect 18556 -2040 19276 -1320
rect 19968 -2040 20688 -1320
rect 21380 -2040 22100 -1320
rect 22792 -2040 23512 -1320
rect -23804 -3160 -23084 -2440
rect -22392 -3160 -21672 -2440
rect -20980 -3160 -20260 -2440
rect -19568 -3160 -18848 -2440
rect -18156 -3160 -17436 -2440
rect -16744 -3160 -16024 -2440
rect -15332 -3160 -14612 -2440
rect -13920 -3160 -13200 -2440
rect -12508 -3160 -11788 -2440
rect -11096 -3160 -10376 -2440
rect -9684 -3160 -8964 -2440
rect -8272 -3160 -7552 -2440
rect -6860 -3160 -6140 -2440
rect -5448 -3160 -4728 -2440
rect -4036 -3160 -3316 -2440
rect -2624 -3160 -1904 -2440
rect -1212 -3160 -492 -2440
rect 200 -3160 920 -2440
rect 1612 -3160 2332 -2440
rect 3024 -3160 3744 -2440
rect 4436 -3160 5156 -2440
rect 5848 -3160 6568 -2440
rect 7260 -3160 7980 -2440
rect 8672 -3160 9392 -2440
rect 10084 -3160 10804 -2440
rect 11496 -3160 12216 -2440
rect 12908 -3160 13628 -2440
rect 14320 -3160 15040 -2440
rect 15732 -3160 16452 -2440
rect 17144 -3160 17864 -2440
rect 18556 -3160 19276 -2440
rect 19968 -3160 20688 -2440
rect 21380 -3160 22100 -2440
rect 22792 -3160 23512 -2440
rect -23804 -4280 -23084 -3560
rect -22392 -4280 -21672 -3560
rect -20980 -4280 -20260 -3560
rect -19568 -4280 -18848 -3560
rect -18156 -4280 -17436 -3560
rect -16744 -4280 -16024 -3560
rect -15332 -4280 -14612 -3560
rect -13920 -4280 -13200 -3560
rect -12508 -4280 -11788 -3560
rect -11096 -4280 -10376 -3560
rect -9684 -4280 -8964 -3560
rect -8272 -4280 -7552 -3560
rect -6860 -4280 -6140 -3560
rect -5448 -4280 -4728 -3560
rect -4036 -4280 -3316 -3560
rect -2624 -4280 -1904 -3560
rect -1212 -4280 -492 -3560
rect 200 -4280 920 -3560
rect 1612 -4280 2332 -3560
rect 3024 -4280 3744 -3560
rect 4436 -4280 5156 -3560
rect 5848 -4280 6568 -3560
rect 7260 -4280 7980 -3560
rect 8672 -4280 9392 -3560
rect 10084 -4280 10804 -3560
rect 11496 -4280 12216 -3560
rect 12908 -4280 13628 -3560
rect 14320 -4280 15040 -3560
rect 15732 -4280 16452 -3560
rect 17144 -4280 17864 -3560
rect 18556 -4280 19276 -3560
rect 19968 -4280 20688 -3560
rect 21380 -4280 22100 -3560
rect 22792 -4280 23512 -3560
rect -23804 -5400 -23084 -4680
rect -22392 -5400 -21672 -4680
rect -20980 -5400 -20260 -4680
rect -19568 -5400 -18848 -4680
rect -18156 -5400 -17436 -4680
rect -16744 -5400 -16024 -4680
rect -15332 -5400 -14612 -4680
rect -13920 -5400 -13200 -4680
rect -12508 -5400 -11788 -4680
rect -11096 -5400 -10376 -4680
rect -9684 -5400 -8964 -4680
rect -8272 -5400 -7552 -4680
rect -6860 -5400 -6140 -4680
rect -5448 -5400 -4728 -4680
rect -4036 -5400 -3316 -4680
rect -2624 -5400 -1904 -4680
rect -1212 -5400 -492 -4680
rect 200 -5400 920 -4680
rect 1612 -5400 2332 -4680
rect 3024 -5400 3744 -4680
rect 4436 -5400 5156 -4680
rect 5848 -5400 6568 -4680
rect 7260 -5400 7980 -4680
rect 8672 -5400 9392 -4680
rect 10084 -5400 10804 -4680
rect 11496 -5400 12216 -4680
rect 12908 -5400 13628 -4680
rect 14320 -5400 15040 -4680
rect 15732 -5400 16452 -4680
rect 17144 -5400 17864 -4680
rect 18556 -5400 19276 -4680
rect 19968 -5400 20688 -4680
rect 21380 -5400 22100 -4680
rect 22792 -5400 23512 -4680
rect -23804 -6520 -23084 -5800
rect -22392 -6520 -21672 -5800
rect -20980 -6520 -20260 -5800
rect -19568 -6520 -18848 -5800
rect -18156 -6520 -17436 -5800
rect -16744 -6520 -16024 -5800
rect -15332 -6520 -14612 -5800
rect -13920 -6520 -13200 -5800
rect -12508 -6520 -11788 -5800
rect -11096 -6520 -10376 -5800
rect -9684 -6520 -8964 -5800
rect -8272 -6520 -7552 -5800
rect -6860 -6520 -6140 -5800
rect -5448 -6520 -4728 -5800
rect -4036 -6520 -3316 -5800
rect -2624 -6520 -1904 -5800
rect -1212 -6520 -492 -5800
rect 200 -6520 920 -5800
rect 1612 -6520 2332 -5800
rect 3024 -6520 3744 -5800
rect 4436 -6520 5156 -5800
rect 5848 -6520 6568 -5800
rect 7260 -6520 7980 -5800
rect 8672 -6520 9392 -5800
rect 10084 -6520 10804 -5800
rect 11496 -6520 12216 -5800
rect 12908 -6520 13628 -5800
rect 14320 -6520 15040 -5800
rect 15732 -6520 16452 -5800
rect 17144 -6520 17864 -5800
rect 18556 -6520 19276 -5800
rect 19968 -6520 20688 -5800
rect 21380 -6520 22100 -5800
rect 22792 -6520 23512 -5800
rect -23804 -7640 -23084 -6920
rect -22392 -7640 -21672 -6920
rect -20980 -7640 -20260 -6920
rect -19568 -7640 -18848 -6920
rect -18156 -7640 -17436 -6920
rect -16744 -7640 -16024 -6920
rect -15332 -7640 -14612 -6920
rect -13920 -7640 -13200 -6920
rect -12508 -7640 -11788 -6920
rect -11096 -7640 -10376 -6920
rect -9684 -7640 -8964 -6920
rect -8272 -7640 -7552 -6920
rect -6860 -7640 -6140 -6920
rect -5448 -7640 -4728 -6920
rect -4036 -7640 -3316 -6920
rect -2624 -7640 -1904 -6920
rect -1212 -7640 -492 -6920
rect 200 -7640 920 -6920
rect 1612 -7640 2332 -6920
rect 3024 -7640 3744 -6920
rect 4436 -7640 5156 -6920
rect 5848 -7640 6568 -6920
rect 7260 -7640 7980 -6920
rect 8672 -7640 9392 -6920
rect 10084 -7640 10804 -6920
rect 11496 -7640 12216 -6920
rect 12908 -7640 13628 -6920
rect 14320 -7640 15040 -6920
rect 15732 -7640 16452 -6920
rect 17144 -7640 17864 -6920
rect 18556 -7640 19276 -6920
rect 19968 -7640 20688 -6920
rect 21380 -7640 22100 -6920
rect 22792 -7640 23512 -6920
rect -23804 -8760 -23084 -8040
rect -22392 -8760 -21672 -8040
rect -20980 -8760 -20260 -8040
rect -19568 -8760 -18848 -8040
rect -18156 -8760 -17436 -8040
rect -16744 -8760 -16024 -8040
rect -15332 -8760 -14612 -8040
rect -13920 -8760 -13200 -8040
rect -12508 -8760 -11788 -8040
rect -11096 -8760 -10376 -8040
rect -9684 -8760 -8964 -8040
rect -8272 -8760 -7552 -8040
rect -6860 -8760 -6140 -8040
rect -5448 -8760 -4728 -8040
rect -4036 -8760 -3316 -8040
rect -2624 -8760 -1904 -8040
rect -1212 -8760 -492 -8040
rect 200 -8760 920 -8040
rect 1612 -8760 2332 -8040
rect 3024 -8760 3744 -8040
rect 4436 -8760 5156 -8040
rect 5848 -8760 6568 -8040
rect 7260 -8760 7980 -8040
rect 8672 -8760 9392 -8040
rect 10084 -8760 10804 -8040
rect 11496 -8760 12216 -8040
rect 12908 -8760 13628 -8040
rect 14320 -8760 15040 -8040
rect 15732 -8760 16452 -8040
rect 17144 -8760 17864 -8040
rect 18556 -8760 19276 -8040
rect 19968 -8760 20688 -8040
rect 21380 -8760 22100 -8040
rect 22792 -8760 23512 -8040
rect -23804 -9880 -23084 -9160
rect -22392 -9880 -21672 -9160
rect -20980 -9880 -20260 -9160
rect -19568 -9880 -18848 -9160
rect -18156 -9880 -17436 -9160
rect -16744 -9880 -16024 -9160
rect -15332 -9880 -14612 -9160
rect -13920 -9880 -13200 -9160
rect -12508 -9880 -11788 -9160
rect -11096 -9880 -10376 -9160
rect -9684 -9880 -8964 -9160
rect -8272 -9880 -7552 -9160
rect -6860 -9880 -6140 -9160
rect -5448 -9880 -4728 -9160
rect -4036 -9880 -3316 -9160
rect -2624 -9880 -1904 -9160
rect -1212 -9880 -492 -9160
rect 200 -9880 920 -9160
rect 1612 -9880 2332 -9160
rect 3024 -9880 3744 -9160
rect 4436 -9880 5156 -9160
rect 5848 -9880 6568 -9160
rect 7260 -9880 7980 -9160
rect 8672 -9880 9392 -9160
rect 10084 -9880 10804 -9160
rect 11496 -9880 12216 -9160
rect 12908 -9880 13628 -9160
rect 14320 -9880 15040 -9160
rect 15732 -9880 16452 -9160
rect 17144 -9880 17864 -9160
rect 18556 -9880 19276 -9160
rect 19968 -9880 20688 -9160
rect 21380 -9880 22100 -9160
rect 22792 -9880 23512 -9160
rect -23804 -11000 -23084 -10280
rect -22392 -11000 -21672 -10280
rect -20980 -11000 -20260 -10280
rect -19568 -11000 -18848 -10280
rect -18156 -11000 -17436 -10280
rect -16744 -11000 -16024 -10280
rect -15332 -11000 -14612 -10280
rect -13920 -11000 -13200 -10280
rect -12508 -11000 -11788 -10280
rect -11096 -11000 -10376 -10280
rect -9684 -11000 -8964 -10280
rect -8272 -11000 -7552 -10280
rect -6860 -11000 -6140 -10280
rect -5448 -11000 -4728 -10280
rect -4036 -11000 -3316 -10280
rect -2624 -11000 -1904 -10280
rect -1212 -11000 -492 -10280
rect 200 -11000 920 -10280
rect 1612 -11000 2332 -10280
rect 3024 -11000 3744 -10280
rect 4436 -11000 5156 -10280
rect 5848 -11000 6568 -10280
rect 7260 -11000 7980 -10280
rect 8672 -11000 9392 -10280
rect 10084 -11000 10804 -10280
rect 11496 -11000 12216 -10280
rect 12908 -11000 13628 -10280
rect 14320 -11000 15040 -10280
rect 15732 -11000 16452 -10280
rect 17144 -11000 17864 -10280
rect 18556 -11000 19276 -10280
rect 19968 -11000 20688 -10280
rect 21380 -11000 22100 -10280
rect 22792 -11000 23512 -10280
rect -23804 -12120 -23084 -11400
rect -22392 -12120 -21672 -11400
rect -20980 -12120 -20260 -11400
rect -19568 -12120 -18848 -11400
rect -18156 -12120 -17436 -11400
rect -16744 -12120 -16024 -11400
rect -15332 -12120 -14612 -11400
rect -13920 -12120 -13200 -11400
rect -12508 -12120 -11788 -11400
rect -11096 -12120 -10376 -11400
rect -9684 -12120 -8964 -11400
rect -8272 -12120 -7552 -11400
rect -6860 -12120 -6140 -11400
rect -5448 -12120 -4728 -11400
rect -4036 -12120 -3316 -11400
rect -2624 -12120 -1904 -11400
rect -1212 -12120 -492 -11400
rect 200 -12120 920 -11400
rect 1612 -12120 2332 -11400
rect 3024 -12120 3744 -11400
rect 4436 -12120 5156 -11400
rect 5848 -12120 6568 -11400
rect 7260 -12120 7980 -11400
rect 8672 -12120 9392 -11400
rect 10084 -12120 10804 -11400
rect 11496 -12120 12216 -11400
rect 12908 -12120 13628 -11400
rect 14320 -12120 15040 -11400
rect 15732 -12120 16452 -11400
rect 17144 -12120 17864 -11400
rect 18556 -12120 19276 -11400
rect 19968 -12120 20688 -11400
rect 21380 -12120 22100 -11400
rect 22792 -12120 23512 -11400
rect -23804 -13240 -23084 -12520
rect -22392 -13240 -21672 -12520
rect -20980 -13240 -20260 -12520
rect -19568 -13240 -18848 -12520
rect -18156 -13240 -17436 -12520
rect -16744 -13240 -16024 -12520
rect -15332 -13240 -14612 -12520
rect -13920 -13240 -13200 -12520
rect -12508 -13240 -11788 -12520
rect -11096 -13240 -10376 -12520
rect -9684 -13240 -8964 -12520
rect -8272 -13240 -7552 -12520
rect -6860 -13240 -6140 -12520
rect -5448 -13240 -4728 -12520
rect -4036 -13240 -3316 -12520
rect -2624 -13240 -1904 -12520
rect -1212 -13240 -492 -12520
rect 200 -13240 920 -12520
rect 1612 -13240 2332 -12520
rect 3024 -13240 3744 -12520
rect 4436 -13240 5156 -12520
rect 5848 -13240 6568 -12520
rect 7260 -13240 7980 -12520
rect 8672 -13240 9392 -12520
rect 10084 -13240 10804 -12520
rect 11496 -13240 12216 -12520
rect 12908 -13240 13628 -12520
rect 14320 -13240 15040 -12520
rect 15732 -13240 16452 -12520
rect 17144 -13240 17864 -12520
rect 18556 -13240 19276 -12520
rect 19968 -13240 20688 -12520
rect 21380 -13240 22100 -12520
rect 22792 -13240 23512 -12520
rect -23804 -14360 -23084 -13640
rect -22392 -14360 -21672 -13640
rect -20980 -14360 -20260 -13640
rect -19568 -14360 -18848 -13640
rect -18156 -14360 -17436 -13640
rect -16744 -14360 -16024 -13640
rect -15332 -14360 -14612 -13640
rect -13920 -14360 -13200 -13640
rect -12508 -14360 -11788 -13640
rect -11096 -14360 -10376 -13640
rect -9684 -14360 -8964 -13640
rect -8272 -14360 -7552 -13640
rect -6860 -14360 -6140 -13640
rect -5448 -14360 -4728 -13640
rect -4036 -14360 -3316 -13640
rect -2624 -14360 -1904 -13640
rect -1212 -14360 -492 -13640
rect 200 -14360 920 -13640
rect 1612 -14360 2332 -13640
rect 3024 -14360 3744 -13640
rect 4436 -14360 5156 -13640
rect 5848 -14360 6568 -13640
rect 7260 -14360 7980 -13640
rect 8672 -14360 9392 -13640
rect 10084 -14360 10804 -13640
rect 11496 -14360 12216 -13640
rect 12908 -14360 13628 -13640
rect 14320 -14360 15040 -13640
rect 15732 -14360 16452 -13640
rect 17144 -14360 17864 -13640
rect 18556 -14360 19276 -13640
rect 19968 -14360 20688 -13640
rect 21380 -14360 22100 -13640
rect 22792 -14360 23512 -13640
rect -23804 -15480 -23084 -14760
rect -22392 -15480 -21672 -14760
rect -20980 -15480 -20260 -14760
rect -19568 -15480 -18848 -14760
rect -18156 -15480 -17436 -14760
rect -16744 -15480 -16024 -14760
rect -15332 -15480 -14612 -14760
rect -13920 -15480 -13200 -14760
rect -12508 -15480 -11788 -14760
rect -11096 -15480 -10376 -14760
rect -9684 -15480 -8964 -14760
rect -8272 -15480 -7552 -14760
rect -6860 -15480 -6140 -14760
rect -5448 -15480 -4728 -14760
rect -4036 -15480 -3316 -14760
rect -2624 -15480 -1904 -14760
rect -1212 -15480 -492 -14760
rect 200 -15480 920 -14760
rect 1612 -15480 2332 -14760
rect 3024 -15480 3744 -14760
rect 4436 -15480 5156 -14760
rect 5848 -15480 6568 -14760
rect 7260 -15480 7980 -14760
rect 8672 -15480 9392 -14760
rect 10084 -15480 10804 -14760
rect 11496 -15480 12216 -14760
rect 12908 -15480 13628 -14760
rect 14320 -15480 15040 -14760
rect 15732 -15480 16452 -14760
rect 17144 -15480 17864 -14760
rect 18556 -15480 19276 -14760
rect 19968 -15480 20688 -14760
rect 21380 -15480 22100 -14760
rect 22792 -15480 23512 -14760
rect -23804 -16600 -23084 -15880
rect -22392 -16600 -21672 -15880
rect -20980 -16600 -20260 -15880
rect -19568 -16600 -18848 -15880
rect -18156 -16600 -17436 -15880
rect -16744 -16600 -16024 -15880
rect -15332 -16600 -14612 -15880
rect -13920 -16600 -13200 -15880
rect -12508 -16600 -11788 -15880
rect -11096 -16600 -10376 -15880
rect -9684 -16600 -8964 -15880
rect -8272 -16600 -7552 -15880
rect -6860 -16600 -6140 -15880
rect -5448 -16600 -4728 -15880
rect -4036 -16600 -3316 -15880
rect -2624 -16600 -1904 -15880
rect -1212 -16600 -492 -15880
rect 200 -16600 920 -15880
rect 1612 -16600 2332 -15880
rect 3024 -16600 3744 -15880
rect 4436 -16600 5156 -15880
rect 5848 -16600 6568 -15880
rect 7260 -16600 7980 -15880
rect 8672 -16600 9392 -15880
rect 10084 -16600 10804 -15880
rect 11496 -16600 12216 -15880
rect 12908 -16600 13628 -15880
rect 14320 -16600 15040 -15880
rect 15732 -16600 16452 -15880
rect 17144 -16600 17864 -15880
rect 18556 -16600 19276 -15880
rect 19968 -16600 20688 -15880
rect 21380 -16600 22100 -15880
rect 22792 -16600 23512 -15880
rect -23804 -17720 -23084 -17000
rect -22392 -17720 -21672 -17000
rect -20980 -17720 -20260 -17000
rect -19568 -17720 -18848 -17000
rect -18156 -17720 -17436 -17000
rect -16744 -17720 -16024 -17000
rect -15332 -17720 -14612 -17000
rect -13920 -17720 -13200 -17000
rect -12508 -17720 -11788 -17000
rect -11096 -17720 -10376 -17000
rect -9684 -17720 -8964 -17000
rect -8272 -17720 -7552 -17000
rect -6860 -17720 -6140 -17000
rect -5448 -17720 -4728 -17000
rect -4036 -17720 -3316 -17000
rect -2624 -17720 -1904 -17000
rect -1212 -17720 -492 -17000
rect 200 -17720 920 -17000
rect 1612 -17720 2332 -17000
rect 3024 -17720 3744 -17000
rect 4436 -17720 5156 -17000
rect 5848 -17720 6568 -17000
rect 7260 -17720 7980 -17000
rect 8672 -17720 9392 -17000
rect 10084 -17720 10804 -17000
rect 11496 -17720 12216 -17000
rect 12908 -17720 13628 -17000
rect 14320 -17720 15040 -17000
rect 15732 -17720 16452 -17000
rect 17144 -17720 17864 -17000
rect 18556 -17720 19276 -17000
rect 19968 -17720 20688 -17000
rect 21380 -17720 22100 -17000
rect 22792 -17720 23512 -17000
rect -23804 -18840 -23084 -18120
rect -22392 -18840 -21672 -18120
rect -20980 -18840 -20260 -18120
rect -19568 -18840 -18848 -18120
rect -18156 -18840 -17436 -18120
rect -16744 -18840 -16024 -18120
rect -15332 -18840 -14612 -18120
rect -13920 -18840 -13200 -18120
rect -12508 -18840 -11788 -18120
rect -11096 -18840 -10376 -18120
rect -9684 -18840 -8964 -18120
rect -8272 -18840 -7552 -18120
rect -6860 -18840 -6140 -18120
rect -5448 -18840 -4728 -18120
rect -4036 -18840 -3316 -18120
rect -2624 -18840 -1904 -18120
rect -1212 -18840 -492 -18120
rect 200 -18840 920 -18120
rect 1612 -18840 2332 -18120
rect 3024 -18840 3744 -18120
rect 4436 -18840 5156 -18120
rect 5848 -18840 6568 -18120
rect 7260 -18840 7980 -18120
rect 8672 -18840 9392 -18120
rect 10084 -18840 10804 -18120
rect 11496 -18840 12216 -18120
rect 12908 -18840 13628 -18120
rect 14320 -18840 15040 -18120
rect 15732 -18840 16452 -18120
rect 17144 -18840 17864 -18120
rect 18556 -18840 19276 -18120
rect 19968 -18840 20688 -18120
rect 21380 -18840 22100 -18120
rect 22792 -18840 23512 -18120
<< metal4 >>
rect -22812 18892 -22716 18908
rect -23805 18840 -23083 18841
rect -23805 18120 -23804 18840
rect -23084 18120 -23083 18840
rect -23805 18119 -23083 18120
rect -22812 18068 -22796 18892
rect -22732 18068 -22716 18892
rect -21400 18892 -21304 18908
rect -22393 18840 -21671 18841
rect -22393 18120 -22392 18840
rect -21672 18120 -21671 18840
rect -22393 18119 -21671 18120
rect -22812 18052 -22716 18068
rect -21400 18068 -21384 18892
rect -21320 18068 -21304 18892
rect -19988 18892 -19892 18908
rect -20981 18840 -20259 18841
rect -20981 18120 -20980 18840
rect -20260 18120 -20259 18840
rect -20981 18119 -20259 18120
rect -21400 18052 -21304 18068
rect -19988 18068 -19972 18892
rect -19908 18068 -19892 18892
rect -18576 18892 -18480 18908
rect -19569 18840 -18847 18841
rect -19569 18120 -19568 18840
rect -18848 18120 -18847 18840
rect -19569 18119 -18847 18120
rect -19988 18052 -19892 18068
rect -18576 18068 -18560 18892
rect -18496 18068 -18480 18892
rect -17164 18892 -17068 18908
rect -18157 18840 -17435 18841
rect -18157 18120 -18156 18840
rect -17436 18120 -17435 18840
rect -18157 18119 -17435 18120
rect -18576 18052 -18480 18068
rect -17164 18068 -17148 18892
rect -17084 18068 -17068 18892
rect -15752 18892 -15656 18908
rect -16745 18840 -16023 18841
rect -16745 18120 -16744 18840
rect -16024 18120 -16023 18840
rect -16745 18119 -16023 18120
rect -17164 18052 -17068 18068
rect -15752 18068 -15736 18892
rect -15672 18068 -15656 18892
rect -14340 18892 -14244 18908
rect -15333 18840 -14611 18841
rect -15333 18120 -15332 18840
rect -14612 18120 -14611 18840
rect -15333 18119 -14611 18120
rect -15752 18052 -15656 18068
rect -14340 18068 -14324 18892
rect -14260 18068 -14244 18892
rect -12928 18892 -12832 18908
rect -13921 18840 -13199 18841
rect -13921 18120 -13920 18840
rect -13200 18120 -13199 18840
rect -13921 18119 -13199 18120
rect -14340 18052 -14244 18068
rect -12928 18068 -12912 18892
rect -12848 18068 -12832 18892
rect -11516 18892 -11420 18908
rect -12509 18840 -11787 18841
rect -12509 18120 -12508 18840
rect -11788 18120 -11787 18840
rect -12509 18119 -11787 18120
rect -12928 18052 -12832 18068
rect -11516 18068 -11500 18892
rect -11436 18068 -11420 18892
rect -10104 18892 -10008 18908
rect -11097 18840 -10375 18841
rect -11097 18120 -11096 18840
rect -10376 18120 -10375 18840
rect -11097 18119 -10375 18120
rect -11516 18052 -11420 18068
rect -10104 18068 -10088 18892
rect -10024 18068 -10008 18892
rect -8692 18892 -8596 18908
rect -9685 18840 -8963 18841
rect -9685 18120 -9684 18840
rect -8964 18120 -8963 18840
rect -9685 18119 -8963 18120
rect -10104 18052 -10008 18068
rect -8692 18068 -8676 18892
rect -8612 18068 -8596 18892
rect -7280 18892 -7184 18908
rect -8273 18840 -7551 18841
rect -8273 18120 -8272 18840
rect -7552 18120 -7551 18840
rect -8273 18119 -7551 18120
rect -8692 18052 -8596 18068
rect -7280 18068 -7264 18892
rect -7200 18068 -7184 18892
rect -5868 18892 -5772 18908
rect -6861 18840 -6139 18841
rect -6861 18120 -6860 18840
rect -6140 18120 -6139 18840
rect -6861 18119 -6139 18120
rect -7280 18052 -7184 18068
rect -5868 18068 -5852 18892
rect -5788 18068 -5772 18892
rect -4456 18892 -4360 18908
rect -5449 18840 -4727 18841
rect -5449 18120 -5448 18840
rect -4728 18120 -4727 18840
rect -5449 18119 -4727 18120
rect -5868 18052 -5772 18068
rect -4456 18068 -4440 18892
rect -4376 18068 -4360 18892
rect -3044 18892 -2948 18908
rect -4037 18840 -3315 18841
rect -4037 18120 -4036 18840
rect -3316 18120 -3315 18840
rect -4037 18119 -3315 18120
rect -4456 18052 -4360 18068
rect -3044 18068 -3028 18892
rect -2964 18068 -2948 18892
rect -1632 18892 -1536 18908
rect -2625 18840 -1903 18841
rect -2625 18120 -2624 18840
rect -1904 18120 -1903 18840
rect -2625 18119 -1903 18120
rect -3044 18052 -2948 18068
rect -1632 18068 -1616 18892
rect -1552 18068 -1536 18892
rect -220 18892 -124 18908
rect -1213 18840 -491 18841
rect -1213 18120 -1212 18840
rect -492 18120 -491 18840
rect -1213 18119 -491 18120
rect -1632 18052 -1536 18068
rect -220 18068 -204 18892
rect -140 18068 -124 18892
rect 1192 18892 1288 18908
rect 199 18840 921 18841
rect 199 18120 200 18840
rect 920 18120 921 18840
rect 199 18119 921 18120
rect -220 18052 -124 18068
rect 1192 18068 1208 18892
rect 1272 18068 1288 18892
rect 2604 18892 2700 18908
rect 1611 18840 2333 18841
rect 1611 18120 1612 18840
rect 2332 18120 2333 18840
rect 1611 18119 2333 18120
rect 1192 18052 1288 18068
rect 2604 18068 2620 18892
rect 2684 18068 2700 18892
rect 4016 18892 4112 18908
rect 3023 18840 3745 18841
rect 3023 18120 3024 18840
rect 3744 18120 3745 18840
rect 3023 18119 3745 18120
rect 2604 18052 2700 18068
rect 4016 18068 4032 18892
rect 4096 18068 4112 18892
rect 5428 18892 5524 18908
rect 4435 18840 5157 18841
rect 4435 18120 4436 18840
rect 5156 18120 5157 18840
rect 4435 18119 5157 18120
rect 4016 18052 4112 18068
rect 5428 18068 5444 18892
rect 5508 18068 5524 18892
rect 6840 18892 6936 18908
rect 5847 18840 6569 18841
rect 5847 18120 5848 18840
rect 6568 18120 6569 18840
rect 5847 18119 6569 18120
rect 5428 18052 5524 18068
rect 6840 18068 6856 18892
rect 6920 18068 6936 18892
rect 8252 18892 8348 18908
rect 7259 18840 7981 18841
rect 7259 18120 7260 18840
rect 7980 18120 7981 18840
rect 7259 18119 7981 18120
rect 6840 18052 6936 18068
rect 8252 18068 8268 18892
rect 8332 18068 8348 18892
rect 9664 18892 9760 18908
rect 8671 18840 9393 18841
rect 8671 18120 8672 18840
rect 9392 18120 9393 18840
rect 8671 18119 9393 18120
rect 8252 18052 8348 18068
rect 9664 18068 9680 18892
rect 9744 18068 9760 18892
rect 11076 18892 11172 18908
rect 10083 18840 10805 18841
rect 10083 18120 10084 18840
rect 10804 18120 10805 18840
rect 10083 18119 10805 18120
rect 9664 18052 9760 18068
rect 11076 18068 11092 18892
rect 11156 18068 11172 18892
rect 12488 18892 12584 18908
rect 11495 18840 12217 18841
rect 11495 18120 11496 18840
rect 12216 18120 12217 18840
rect 11495 18119 12217 18120
rect 11076 18052 11172 18068
rect 12488 18068 12504 18892
rect 12568 18068 12584 18892
rect 13900 18892 13996 18908
rect 12907 18840 13629 18841
rect 12907 18120 12908 18840
rect 13628 18120 13629 18840
rect 12907 18119 13629 18120
rect 12488 18052 12584 18068
rect 13900 18068 13916 18892
rect 13980 18068 13996 18892
rect 15312 18892 15408 18908
rect 14319 18840 15041 18841
rect 14319 18120 14320 18840
rect 15040 18120 15041 18840
rect 14319 18119 15041 18120
rect 13900 18052 13996 18068
rect 15312 18068 15328 18892
rect 15392 18068 15408 18892
rect 16724 18892 16820 18908
rect 15731 18840 16453 18841
rect 15731 18120 15732 18840
rect 16452 18120 16453 18840
rect 15731 18119 16453 18120
rect 15312 18052 15408 18068
rect 16724 18068 16740 18892
rect 16804 18068 16820 18892
rect 18136 18892 18232 18908
rect 17143 18840 17865 18841
rect 17143 18120 17144 18840
rect 17864 18120 17865 18840
rect 17143 18119 17865 18120
rect 16724 18052 16820 18068
rect 18136 18068 18152 18892
rect 18216 18068 18232 18892
rect 19548 18892 19644 18908
rect 18555 18840 19277 18841
rect 18555 18120 18556 18840
rect 19276 18120 19277 18840
rect 18555 18119 19277 18120
rect 18136 18052 18232 18068
rect 19548 18068 19564 18892
rect 19628 18068 19644 18892
rect 20960 18892 21056 18908
rect 19967 18840 20689 18841
rect 19967 18120 19968 18840
rect 20688 18120 20689 18840
rect 19967 18119 20689 18120
rect 19548 18052 19644 18068
rect 20960 18068 20976 18892
rect 21040 18068 21056 18892
rect 22372 18892 22468 18908
rect 21379 18840 22101 18841
rect 21379 18120 21380 18840
rect 22100 18120 22101 18840
rect 21379 18119 22101 18120
rect 20960 18052 21056 18068
rect 22372 18068 22388 18892
rect 22452 18068 22468 18892
rect 23784 18892 23880 18908
rect 22791 18840 23513 18841
rect 22791 18120 22792 18840
rect 23512 18120 23513 18840
rect 22791 18119 23513 18120
rect 22372 18052 22468 18068
rect 23784 18068 23800 18892
rect 23864 18068 23880 18892
rect 23784 18052 23880 18068
rect -22812 17772 -22716 17788
rect -23805 17720 -23083 17721
rect -23805 17000 -23804 17720
rect -23084 17000 -23083 17720
rect -23805 16999 -23083 17000
rect -22812 16948 -22796 17772
rect -22732 16948 -22716 17772
rect -21400 17772 -21304 17788
rect -22393 17720 -21671 17721
rect -22393 17000 -22392 17720
rect -21672 17000 -21671 17720
rect -22393 16999 -21671 17000
rect -22812 16932 -22716 16948
rect -21400 16948 -21384 17772
rect -21320 16948 -21304 17772
rect -19988 17772 -19892 17788
rect -20981 17720 -20259 17721
rect -20981 17000 -20980 17720
rect -20260 17000 -20259 17720
rect -20981 16999 -20259 17000
rect -21400 16932 -21304 16948
rect -19988 16948 -19972 17772
rect -19908 16948 -19892 17772
rect -18576 17772 -18480 17788
rect -19569 17720 -18847 17721
rect -19569 17000 -19568 17720
rect -18848 17000 -18847 17720
rect -19569 16999 -18847 17000
rect -19988 16932 -19892 16948
rect -18576 16948 -18560 17772
rect -18496 16948 -18480 17772
rect -17164 17772 -17068 17788
rect -18157 17720 -17435 17721
rect -18157 17000 -18156 17720
rect -17436 17000 -17435 17720
rect -18157 16999 -17435 17000
rect -18576 16932 -18480 16948
rect -17164 16948 -17148 17772
rect -17084 16948 -17068 17772
rect -15752 17772 -15656 17788
rect -16745 17720 -16023 17721
rect -16745 17000 -16744 17720
rect -16024 17000 -16023 17720
rect -16745 16999 -16023 17000
rect -17164 16932 -17068 16948
rect -15752 16948 -15736 17772
rect -15672 16948 -15656 17772
rect -14340 17772 -14244 17788
rect -15333 17720 -14611 17721
rect -15333 17000 -15332 17720
rect -14612 17000 -14611 17720
rect -15333 16999 -14611 17000
rect -15752 16932 -15656 16948
rect -14340 16948 -14324 17772
rect -14260 16948 -14244 17772
rect -12928 17772 -12832 17788
rect -13921 17720 -13199 17721
rect -13921 17000 -13920 17720
rect -13200 17000 -13199 17720
rect -13921 16999 -13199 17000
rect -14340 16932 -14244 16948
rect -12928 16948 -12912 17772
rect -12848 16948 -12832 17772
rect -11516 17772 -11420 17788
rect -12509 17720 -11787 17721
rect -12509 17000 -12508 17720
rect -11788 17000 -11787 17720
rect -12509 16999 -11787 17000
rect -12928 16932 -12832 16948
rect -11516 16948 -11500 17772
rect -11436 16948 -11420 17772
rect -10104 17772 -10008 17788
rect -11097 17720 -10375 17721
rect -11097 17000 -11096 17720
rect -10376 17000 -10375 17720
rect -11097 16999 -10375 17000
rect -11516 16932 -11420 16948
rect -10104 16948 -10088 17772
rect -10024 16948 -10008 17772
rect -8692 17772 -8596 17788
rect -9685 17720 -8963 17721
rect -9685 17000 -9684 17720
rect -8964 17000 -8963 17720
rect -9685 16999 -8963 17000
rect -10104 16932 -10008 16948
rect -8692 16948 -8676 17772
rect -8612 16948 -8596 17772
rect -7280 17772 -7184 17788
rect -8273 17720 -7551 17721
rect -8273 17000 -8272 17720
rect -7552 17000 -7551 17720
rect -8273 16999 -7551 17000
rect -8692 16932 -8596 16948
rect -7280 16948 -7264 17772
rect -7200 16948 -7184 17772
rect -5868 17772 -5772 17788
rect -6861 17720 -6139 17721
rect -6861 17000 -6860 17720
rect -6140 17000 -6139 17720
rect -6861 16999 -6139 17000
rect -7280 16932 -7184 16948
rect -5868 16948 -5852 17772
rect -5788 16948 -5772 17772
rect -4456 17772 -4360 17788
rect -5449 17720 -4727 17721
rect -5449 17000 -5448 17720
rect -4728 17000 -4727 17720
rect -5449 16999 -4727 17000
rect -5868 16932 -5772 16948
rect -4456 16948 -4440 17772
rect -4376 16948 -4360 17772
rect -3044 17772 -2948 17788
rect -4037 17720 -3315 17721
rect -4037 17000 -4036 17720
rect -3316 17000 -3315 17720
rect -4037 16999 -3315 17000
rect -4456 16932 -4360 16948
rect -3044 16948 -3028 17772
rect -2964 16948 -2948 17772
rect -1632 17772 -1536 17788
rect -2625 17720 -1903 17721
rect -2625 17000 -2624 17720
rect -1904 17000 -1903 17720
rect -2625 16999 -1903 17000
rect -3044 16932 -2948 16948
rect -1632 16948 -1616 17772
rect -1552 16948 -1536 17772
rect -220 17772 -124 17788
rect -1213 17720 -491 17721
rect -1213 17000 -1212 17720
rect -492 17000 -491 17720
rect -1213 16999 -491 17000
rect -1632 16932 -1536 16948
rect -220 16948 -204 17772
rect -140 16948 -124 17772
rect 1192 17772 1288 17788
rect 199 17720 921 17721
rect 199 17000 200 17720
rect 920 17000 921 17720
rect 199 16999 921 17000
rect -220 16932 -124 16948
rect 1192 16948 1208 17772
rect 1272 16948 1288 17772
rect 2604 17772 2700 17788
rect 1611 17720 2333 17721
rect 1611 17000 1612 17720
rect 2332 17000 2333 17720
rect 1611 16999 2333 17000
rect 1192 16932 1288 16948
rect 2604 16948 2620 17772
rect 2684 16948 2700 17772
rect 4016 17772 4112 17788
rect 3023 17720 3745 17721
rect 3023 17000 3024 17720
rect 3744 17000 3745 17720
rect 3023 16999 3745 17000
rect 2604 16932 2700 16948
rect 4016 16948 4032 17772
rect 4096 16948 4112 17772
rect 5428 17772 5524 17788
rect 4435 17720 5157 17721
rect 4435 17000 4436 17720
rect 5156 17000 5157 17720
rect 4435 16999 5157 17000
rect 4016 16932 4112 16948
rect 5428 16948 5444 17772
rect 5508 16948 5524 17772
rect 6840 17772 6936 17788
rect 5847 17720 6569 17721
rect 5847 17000 5848 17720
rect 6568 17000 6569 17720
rect 5847 16999 6569 17000
rect 5428 16932 5524 16948
rect 6840 16948 6856 17772
rect 6920 16948 6936 17772
rect 8252 17772 8348 17788
rect 7259 17720 7981 17721
rect 7259 17000 7260 17720
rect 7980 17000 7981 17720
rect 7259 16999 7981 17000
rect 6840 16932 6936 16948
rect 8252 16948 8268 17772
rect 8332 16948 8348 17772
rect 9664 17772 9760 17788
rect 8671 17720 9393 17721
rect 8671 17000 8672 17720
rect 9392 17000 9393 17720
rect 8671 16999 9393 17000
rect 8252 16932 8348 16948
rect 9664 16948 9680 17772
rect 9744 16948 9760 17772
rect 11076 17772 11172 17788
rect 10083 17720 10805 17721
rect 10083 17000 10084 17720
rect 10804 17000 10805 17720
rect 10083 16999 10805 17000
rect 9664 16932 9760 16948
rect 11076 16948 11092 17772
rect 11156 16948 11172 17772
rect 12488 17772 12584 17788
rect 11495 17720 12217 17721
rect 11495 17000 11496 17720
rect 12216 17000 12217 17720
rect 11495 16999 12217 17000
rect 11076 16932 11172 16948
rect 12488 16948 12504 17772
rect 12568 16948 12584 17772
rect 13900 17772 13996 17788
rect 12907 17720 13629 17721
rect 12907 17000 12908 17720
rect 13628 17000 13629 17720
rect 12907 16999 13629 17000
rect 12488 16932 12584 16948
rect 13900 16948 13916 17772
rect 13980 16948 13996 17772
rect 15312 17772 15408 17788
rect 14319 17720 15041 17721
rect 14319 17000 14320 17720
rect 15040 17000 15041 17720
rect 14319 16999 15041 17000
rect 13900 16932 13996 16948
rect 15312 16948 15328 17772
rect 15392 16948 15408 17772
rect 16724 17772 16820 17788
rect 15731 17720 16453 17721
rect 15731 17000 15732 17720
rect 16452 17000 16453 17720
rect 15731 16999 16453 17000
rect 15312 16932 15408 16948
rect 16724 16948 16740 17772
rect 16804 16948 16820 17772
rect 18136 17772 18232 17788
rect 17143 17720 17865 17721
rect 17143 17000 17144 17720
rect 17864 17000 17865 17720
rect 17143 16999 17865 17000
rect 16724 16932 16820 16948
rect 18136 16948 18152 17772
rect 18216 16948 18232 17772
rect 19548 17772 19644 17788
rect 18555 17720 19277 17721
rect 18555 17000 18556 17720
rect 19276 17000 19277 17720
rect 18555 16999 19277 17000
rect 18136 16932 18232 16948
rect 19548 16948 19564 17772
rect 19628 16948 19644 17772
rect 20960 17772 21056 17788
rect 19967 17720 20689 17721
rect 19967 17000 19968 17720
rect 20688 17000 20689 17720
rect 19967 16999 20689 17000
rect 19548 16932 19644 16948
rect 20960 16948 20976 17772
rect 21040 16948 21056 17772
rect 22372 17772 22468 17788
rect 21379 17720 22101 17721
rect 21379 17000 21380 17720
rect 22100 17000 22101 17720
rect 21379 16999 22101 17000
rect 20960 16932 21056 16948
rect 22372 16948 22388 17772
rect 22452 16948 22468 17772
rect 23784 17772 23880 17788
rect 22791 17720 23513 17721
rect 22791 17000 22792 17720
rect 23512 17000 23513 17720
rect 22791 16999 23513 17000
rect 22372 16932 22468 16948
rect 23784 16948 23800 17772
rect 23864 16948 23880 17772
rect 23784 16932 23880 16948
rect -22812 16652 -22716 16668
rect -23805 16600 -23083 16601
rect -23805 15880 -23804 16600
rect -23084 15880 -23083 16600
rect -23805 15879 -23083 15880
rect -22812 15828 -22796 16652
rect -22732 15828 -22716 16652
rect -21400 16652 -21304 16668
rect -22393 16600 -21671 16601
rect -22393 15880 -22392 16600
rect -21672 15880 -21671 16600
rect -22393 15879 -21671 15880
rect -22812 15812 -22716 15828
rect -21400 15828 -21384 16652
rect -21320 15828 -21304 16652
rect -19988 16652 -19892 16668
rect -20981 16600 -20259 16601
rect -20981 15880 -20980 16600
rect -20260 15880 -20259 16600
rect -20981 15879 -20259 15880
rect -21400 15812 -21304 15828
rect -19988 15828 -19972 16652
rect -19908 15828 -19892 16652
rect -18576 16652 -18480 16668
rect -19569 16600 -18847 16601
rect -19569 15880 -19568 16600
rect -18848 15880 -18847 16600
rect -19569 15879 -18847 15880
rect -19988 15812 -19892 15828
rect -18576 15828 -18560 16652
rect -18496 15828 -18480 16652
rect -17164 16652 -17068 16668
rect -18157 16600 -17435 16601
rect -18157 15880 -18156 16600
rect -17436 15880 -17435 16600
rect -18157 15879 -17435 15880
rect -18576 15812 -18480 15828
rect -17164 15828 -17148 16652
rect -17084 15828 -17068 16652
rect -15752 16652 -15656 16668
rect -16745 16600 -16023 16601
rect -16745 15880 -16744 16600
rect -16024 15880 -16023 16600
rect -16745 15879 -16023 15880
rect -17164 15812 -17068 15828
rect -15752 15828 -15736 16652
rect -15672 15828 -15656 16652
rect -14340 16652 -14244 16668
rect -15333 16600 -14611 16601
rect -15333 15880 -15332 16600
rect -14612 15880 -14611 16600
rect -15333 15879 -14611 15880
rect -15752 15812 -15656 15828
rect -14340 15828 -14324 16652
rect -14260 15828 -14244 16652
rect -12928 16652 -12832 16668
rect -13921 16600 -13199 16601
rect -13921 15880 -13920 16600
rect -13200 15880 -13199 16600
rect -13921 15879 -13199 15880
rect -14340 15812 -14244 15828
rect -12928 15828 -12912 16652
rect -12848 15828 -12832 16652
rect -11516 16652 -11420 16668
rect -12509 16600 -11787 16601
rect -12509 15880 -12508 16600
rect -11788 15880 -11787 16600
rect -12509 15879 -11787 15880
rect -12928 15812 -12832 15828
rect -11516 15828 -11500 16652
rect -11436 15828 -11420 16652
rect -10104 16652 -10008 16668
rect -11097 16600 -10375 16601
rect -11097 15880 -11096 16600
rect -10376 15880 -10375 16600
rect -11097 15879 -10375 15880
rect -11516 15812 -11420 15828
rect -10104 15828 -10088 16652
rect -10024 15828 -10008 16652
rect -8692 16652 -8596 16668
rect -9685 16600 -8963 16601
rect -9685 15880 -9684 16600
rect -8964 15880 -8963 16600
rect -9685 15879 -8963 15880
rect -10104 15812 -10008 15828
rect -8692 15828 -8676 16652
rect -8612 15828 -8596 16652
rect -7280 16652 -7184 16668
rect -8273 16600 -7551 16601
rect -8273 15880 -8272 16600
rect -7552 15880 -7551 16600
rect -8273 15879 -7551 15880
rect -8692 15812 -8596 15828
rect -7280 15828 -7264 16652
rect -7200 15828 -7184 16652
rect -5868 16652 -5772 16668
rect -6861 16600 -6139 16601
rect -6861 15880 -6860 16600
rect -6140 15880 -6139 16600
rect -6861 15879 -6139 15880
rect -7280 15812 -7184 15828
rect -5868 15828 -5852 16652
rect -5788 15828 -5772 16652
rect -4456 16652 -4360 16668
rect -5449 16600 -4727 16601
rect -5449 15880 -5448 16600
rect -4728 15880 -4727 16600
rect -5449 15879 -4727 15880
rect -5868 15812 -5772 15828
rect -4456 15828 -4440 16652
rect -4376 15828 -4360 16652
rect -3044 16652 -2948 16668
rect -4037 16600 -3315 16601
rect -4037 15880 -4036 16600
rect -3316 15880 -3315 16600
rect -4037 15879 -3315 15880
rect -4456 15812 -4360 15828
rect -3044 15828 -3028 16652
rect -2964 15828 -2948 16652
rect -1632 16652 -1536 16668
rect -2625 16600 -1903 16601
rect -2625 15880 -2624 16600
rect -1904 15880 -1903 16600
rect -2625 15879 -1903 15880
rect -3044 15812 -2948 15828
rect -1632 15828 -1616 16652
rect -1552 15828 -1536 16652
rect -220 16652 -124 16668
rect -1213 16600 -491 16601
rect -1213 15880 -1212 16600
rect -492 15880 -491 16600
rect -1213 15879 -491 15880
rect -1632 15812 -1536 15828
rect -220 15828 -204 16652
rect -140 15828 -124 16652
rect 1192 16652 1288 16668
rect 199 16600 921 16601
rect 199 15880 200 16600
rect 920 15880 921 16600
rect 199 15879 921 15880
rect -220 15812 -124 15828
rect 1192 15828 1208 16652
rect 1272 15828 1288 16652
rect 2604 16652 2700 16668
rect 1611 16600 2333 16601
rect 1611 15880 1612 16600
rect 2332 15880 2333 16600
rect 1611 15879 2333 15880
rect 1192 15812 1288 15828
rect 2604 15828 2620 16652
rect 2684 15828 2700 16652
rect 4016 16652 4112 16668
rect 3023 16600 3745 16601
rect 3023 15880 3024 16600
rect 3744 15880 3745 16600
rect 3023 15879 3745 15880
rect 2604 15812 2700 15828
rect 4016 15828 4032 16652
rect 4096 15828 4112 16652
rect 5428 16652 5524 16668
rect 4435 16600 5157 16601
rect 4435 15880 4436 16600
rect 5156 15880 5157 16600
rect 4435 15879 5157 15880
rect 4016 15812 4112 15828
rect 5428 15828 5444 16652
rect 5508 15828 5524 16652
rect 6840 16652 6936 16668
rect 5847 16600 6569 16601
rect 5847 15880 5848 16600
rect 6568 15880 6569 16600
rect 5847 15879 6569 15880
rect 5428 15812 5524 15828
rect 6840 15828 6856 16652
rect 6920 15828 6936 16652
rect 8252 16652 8348 16668
rect 7259 16600 7981 16601
rect 7259 15880 7260 16600
rect 7980 15880 7981 16600
rect 7259 15879 7981 15880
rect 6840 15812 6936 15828
rect 8252 15828 8268 16652
rect 8332 15828 8348 16652
rect 9664 16652 9760 16668
rect 8671 16600 9393 16601
rect 8671 15880 8672 16600
rect 9392 15880 9393 16600
rect 8671 15879 9393 15880
rect 8252 15812 8348 15828
rect 9664 15828 9680 16652
rect 9744 15828 9760 16652
rect 11076 16652 11172 16668
rect 10083 16600 10805 16601
rect 10083 15880 10084 16600
rect 10804 15880 10805 16600
rect 10083 15879 10805 15880
rect 9664 15812 9760 15828
rect 11076 15828 11092 16652
rect 11156 15828 11172 16652
rect 12488 16652 12584 16668
rect 11495 16600 12217 16601
rect 11495 15880 11496 16600
rect 12216 15880 12217 16600
rect 11495 15879 12217 15880
rect 11076 15812 11172 15828
rect 12488 15828 12504 16652
rect 12568 15828 12584 16652
rect 13900 16652 13996 16668
rect 12907 16600 13629 16601
rect 12907 15880 12908 16600
rect 13628 15880 13629 16600
rect 12907 15879 13629 15880
rect 12488 15812 12584 15828
rect 13900 15828 13916 16652
rect 13980 15828 13996 16652
rect 15312 16652 15408 16668
rect 14319 16600 15041 16601
rect 14319 15880 14320 16600
rect 15040 15880 15041 16600
rect 14319 15879 15041 15880
rect 13900 15812 13996 15828
rect 15312 15828 15328 16652
rect 15392 15828 15408 16652
rect 16724 16652 16820 16668
rect 15731 16600 16453 16601
rect 15731 15880 15732 16600
rect 16452 15880 16453 16600
rect 15731 15879 16453 15880
rect 15312 15812 15408 15828
rect 16724 15828 16740 16652
rect 16804 15828 16820 16652
rect 18136 16652 18232 16668
rect 17143 16600 17865 16601
rect 17143 15880 17144 16600
rect 17864 15880 17865 16600
rect 17143 15879 17865 15880
rect 16724 15812 16820 15828
rect 18136 15828 18152 16652
rect 18216 15828 18232 16652
rect 19548 16652 19644 16668
rect 18555 16600 19277 16601
rect 18555 15880 18556 16600
rect 19276 15880 19277 16600
rect 18555 15879 19277 15880
rect 18136 15812 18232 15828
rect 19548 15828 19564 16652
rect 19628 15828 19644 16652
rect 20960 16652 21056 16668
rect 19967 16600 20689 16601
rect 19967 15880 19968 16600
rect 20688 15880 20689 16600
rect 19967 15879 20689 15880
rect 19548 15812 19644 15828
rect 20960 15828 20976 16652
rect 21040 15828 21056 16652
rect 22372 16652 22468 16668
rect 21379 16600 22101 16601
rect 21379 15880 21380 16600
rect 22100 15880 22101 16600
rect 21379 15879 22101 15880
rect 20960 15812 21056 15828
rect 22372 15828 22388 16652
rect 22452 15828 22468 16652
rect 23784 16652 23880 16668
rect 22791 16600 23513 16601
rect 22791 15880 22792 16600
rect 23512 15880 23513 16600
rect 22791 15879 23513 15880
rect 22372 15812 22468 15828
rect 23784 15828 23800 16652
rect 23864 15828 23880 16652
rect 23784 15812 23880 15828
rect -22812 15532 -22716 15548
rect -23805 15480 -23083 15481
rect -23805 14760 -23804 15480
rect -23084 14760 -23083 15480
rect -23805 14759 -23083 14760
rect -22812 14708 -22796 15532
rect -22732 14708 -22716 15532
rect -21400 15532 -21304 15548
rect -22393 15480 -21671 15481
rect -22393 14760 -22392 15480
rect -21672 14760 -21671 15480
rect -22393 14759 -21671 14760
rect -22812 14692 -22716 14708
rect -21400 14708 -21384 15532
rect -21320 14708 -21304 15532
rect -19988 15532 -19892 15548
rect -20981 15480 -20259 15481
rect -20981 14760 -20980 15480
rect -20260 14760 -20259 15480
rect -20981 14759 -20259 14760
rect -21400 14692 -21304 14708
rect -19988 14708 -19972 15532
rect -19908 14708 -19892 15532
rect -18576 15532 -18480 15548
rect -19569 15480 -18847 15481
rect -19569 14760 -19568 15480
rect -18848 14760 -18847 15480
rect -19569 14759 -18847 14760
rect -19988 14692 -19892 14708
rect -18576 14708 -18560 15532
rect -18496 14708 -18480 15532
rect -17164 15532 -17068 15548
rect -18157 15480 -17435 15481
rect -18157 14760 -18156 15480
rect -17436 14760 -17435 15480
rect -18157 14759 -17435 14760
rect -18576 14692 -18480 14708
rect -17164 14708 -17148 15532
rect -17084 14708 -17068 15532
rect -15752 15532 -15656 15548
rect -16745 15480 -16023 15481
rect -16745 14760 -16744 15480
rect -16024 14760 -16023 15480
rect -16745 14759 -16023 14760
rect -17164 14692 -17068 14708
rect -15752 14708 -15736 15532
rect -15672 14708 -15656 15532
rect -14340 15532 -14244 15548
rect -15333 15480 -14611 15481
rect -15333 14760 -15332 15480
rect -14612 14760 -14611 15480
rect -15333 14759 -14611 14760
rect -15752 14692 -15656 14708
rect -14340 14708 -14324 15532
rect -14260 14708 -14244 15532
rect -12928 15532 -12832 15548
rect -13921 15480 -13199 15481
rect -13921 14760 -13920 15480
rect -13200 14760 -13199 15480
rect -13921 14759 -13199 14760
rect -14340 14692 -14244 14708
rect -12928 14708 -12912 15532
rect -12848 14708 -12832 15532
rect -11516 15532 -11420 15548
rect -12509 15480 -11787 15481
rect -12509 14760 -12508 15480
rect -11788 14760 -11787 15480
rect -12509 14759 -11787 14760
rect -12928 14692 -12832 14708
rect -11516 14708 -11500 15532
rect -11436 14708 -11420 15532
rect -10104 15532 -10008 15548
rect -11097 15480 -10375 15481
rect -11097 14760 -11096 15480
rect -10376 14760 -10375 15480
rect -11097 14759 -10375 14760
rect -11516 14692 -11420 14708
rect -10104 14708 -10088 15532
rect -10024 14708 -10008 15532
rect -8692 15532 -8596 15548
rect -9685 15480 -8963 15481
rect -9685 14760 -9684 15480
rect -8964 14760 -8963 15480
rect -9685 14759 -8963 14760
rect -10104 14692 -10008 14708
rect -8692 14708 -8676 15532
rect -8612 14708 -8596 15532
rect -7280 15532 -7184 15548
rect -8273 15480 -7551 15481
rect -8273 14760 -8272 15480
rect -7552 14760 -7551 15480
rect -8273 14759 -7551 14760
rect -8692 14692 -8596 14708
rect -7280 14708 -7264 15532
rect -7200 14708 -7184 15532
rect -5868 15532 -5772 15548
rect -6861 15480 -6139 15481
rect -6861 14760 -6860 15480
rect -6140 14760 -6139 15480
rect -6861 14759 -6139 14760
rect -7280 14692 -7184 14708
rect -5868 14708 -5852 15532
rect -5788 14708 -5772 15532
rect -4456 15532 -4360 15548
rect -5449 15480 -4727 15481
rect -5449 14760 -5448 15480
rect -4728 14760 -4727 15480
rect -5449 14759 -4727 14760
rect -5868 14692 -5772 14708
rect -4456 14708 -4440 15532
rect -4376 14708 -4360 15532
rect -3044 15532 -2948 15548
rect -4037 15480 -3315 15481
rect -4037 14760 -4036 15480
rect -3316 14760 -3315 15480
rect -4037 14759 -3315 14760
rect -4456 14692 -4360 14708
rect -3044 14708 -3028 15532
rect -2964 14708 -2948 15532
rect -1632 15532 -1536 15548
rect -2625 15480 -1903 15481
rect -2625 14760 -2624 15480
rect -1904 14760 -1903 15480
rect -2625 14759 -1903 14760
rect -3044 14692 -2948 14708
rect -1632 14708 -1616 15532
rect -1552 14708 -1536 15532
rect -220 15532 -124 15548
rect -1213 15480 -491 15481
rect -1213 14760 -1212 15480
rect -492 14760 -491 15480
rect -1213 14759 -491 14760
rect -1632 14692 -1536 14708
rect -220 14708 -204 15532
rect -140 14708 -124 15532
rect 1192 15532 1288 15548
rect 199 15480 921 15481
rect 199 14760 200 15480
rect 920 14760 921 15480
rect 199 14759 921 14760
rect -220 14692 -124 14708
rect 1192 14708 1208 15532
rect 1272 14708 1288 15532
rect 2604 15532 2700 15548
rect 1611 15480 2333 15481
rect 1611 14760 1612 15480
rect 2332 14760 2333 15480
rect 1611 14759 2333 14760
rect 1192 14692 1288 14708
rect 2604 14708 2620 15532
rect 2684 14708 2700 15532
rect 4016 15532 4112 15548
rect 3023 15480 3745 15481
rect 3023 14760 3024 15480
rect 3744 14760 3745 15480
rect 3023 14759 3745 14760
rect 2604 14692 2700 14708
rect 4016 14708 4032 15532
rect 4096 14708 4112 15532
rect 5428 15532 5524 15548
rect 4435 15480 5157 15481
rect 4435 14760 4436 15480
rect 5156 14760 5157 15480
rect 4435 14759 5157 14760
rect 4016 14692 4112 14708
rect 5428 14708 5444 15532
rect 5508 14708 5524 15532
rect 6840 15532 6936 15548
rect 5847 15480 6569 15481
rect 5847 14760 5848 15480
rect 6568 14760 6569 15480
rect 5847 14759 6569 14760
rect 5428 14692 5524 14708
rect 6840 14708 6856 15532
rect 6920 14708 6936 15532
rect 8252 15532 8348 15548
rect 7259 15480 7981 15481
rect 7259 14760 7260 15480
rect 7980 14760 7981 15480
rect 7259 14759 7981 14760
rect 6840 14692 6936 14708
rect 8252 14708 8268 15532
rect 8332 14708 8348 15532
rect 9664 15532 9760 15548
rect 8671 15480 9393 15481
rect 8671 14760 8672 15480
rect 9392 14760 9393 15480
rect 8671 14759 9393 14760
rect 8252 14692 8348 14708
rect 9664 14708 9680 15532
rect 9744 14708 9760 15532
rect 11076 15532 11172 15548
rect 10083 15480 10805 15481
rect 10083 14760 10084 15480
rect 10804 14760 10805 15480
rect 10083 14759 10805 14760
rect 9664 14692 9760 14708
rect 11076 14708 11092 15532
rect 11156 14708 11172 15532
rect 12488 15532 12584 15548
rect 11495 15480 12217 15481
rect 11495 14760 11496 15480
rect 12216 14760 12217 15480
rect 11495 14759 12217 14760
rect 11076 14692 11172 14708
rect 12488 14708 12504 15532
rect 12568 14708 12584 15532
rect 13900 15532 13996 15548
rect 12907 15480 13629 15481
rect 12907 14760 12908 15480
rect 13628 14760 13629 15480
rect 12907 14759 13629 14760
rect 12488 14692 12584 14708
rect 13900 14708 13916 15532
rect 13980 14708 13996 15532
rect 15312 15532 15408 15548
rect 14319 15480 15041 15481
rect 14319 14760 14320 15480
rect 15040 14760 15041 15480
rect 14319 14759 15041 14760
rect 13900 14692 13996 14708
rect 15312 14708 15328 15532
rect 15392 14708 15408 15532
rect 16724 15532 16820 15548
rect 15731 15480 16453 15481
rect 15731 14760 15732 15480
rect 16452 14760 16453 15480
rect 15731 14759 16453 14760
rect 15312 14692 15408 14708
rect 16724 14708 16740 15532
rect 16804 14708 16820 15532
rect 18136 15532 18232 15548
rect 17143 15480 17865 15481
rect 17143 14760 17144 15480
rect 17864 14760 17865 15480
rect 17143 14759 17865 14760
rect 16724 14692 16820 14708
rect 18136 14708 18152 15532
rect 18216 14708 18232 15532
rect 19548 15532 19644 15548
rect 18555 15480 19277 15481
rect 18555 14760 18556 15480
rect 19276 14760 19277 15480
rect 18555 14759 19277 14760
rect 18136 14692 18232 14708
rect 19548 14708 19564 15532
rect 19628 14708 19644 15532
rect 20960 15532 21056 15548
rect 19967 15480 20689 15481
rect 19967 14760 19968 15480
rect 20688 14760 20689 15480
rect 19967 14759 20689 14760
rect 19548 14692 19644 14708
rect 20960 14708 20976 15532
rect 21040 14708 21056 15532
rect 22372 15532 22468 15548
rect 21379 15480 22101 15481
rect 21379 14760 21380 15480
rect 22100 14760 22101 15480
rect 21379 14759 22101 14760
rect 20960 14692 21056 14708
rect 22372 14708 22388 15532
rect 22452 14708 22468 15532
rect 23784 15532 23880 15548
rect 22791 15480 23513 15481
rect 22791 14760 22792 15480
rect 23512 14760 23513 15480
rect 22791 14759 23513 14760
rect 22372 14692 22468 14708
rect 23784 14708 23800 15532
rect 23864 14708 23880 15532
rect 23784 14692 23880 14708
rect -22812 14412 -22716 14428
rect -23805 14360 -23083 14361
rect -23805 13640 -23804 14360
rect -23084 13640 -23083 14360
rect -23805 13639 -23083 13640
rect -22812 13588 -22796 14412
rect -22732 13588 -22716 14412
rect -21400 14412 -21304 14428
rect -22393 14360 -21671 14361
rect -22393 13640 -22392 14360
rect -21672 13640 -21671 14360
rect -22393 13639 -21671 13640
rect -22812 13572 -22716 13588
rect -21400 13588 -21384 14412
rect -21320 13588 -21304 14412
rect -19988 14412 -19892 14428
rect -20981 14360 -20259 14361
rect -20981 13640 -20980 14360
rect -20260 13640 -20259 14360
rect -20981 13639 -20259 13640
rect -21400 13572 -21304 13588
rect -19988 13588 -19972 14412
rect -19908 13588 -19892 14412
rect -18576 14412 -18480 14428
rect -19569 14360 -18847 14361
rect -19569 13640 -19568 14360
rect -18848 13640 -18847 14360
rect -19569 13639 -18847 13640
rect -19988 13572 -19892 13588
rect -18576 13588 -18560 14412
rect -18496 13588 -18480 14412
rect -17164 14412 -17068 14428
rect -18157 14360 -17435 14361
rect -18157 13640 -18156 14360
rect -17436 13640 -17435 14360
rect -18157 13639 -17435 13640
rect -18576 13572 -18480 13588
rect -17164 13588 -17148 14412
rect -17084 13588 -17068 14412
rect -15752 14412 -15656 14428
rect -16745 14360 -16023 14361
rect -16745 13640 -16744 14360
rect -16024 13640 -16023 14360
rect -16745 13639 -16023 13640
rect -17164 13572 -17068 13588
rect -15752 13588 -15736 14412
rect -15672 13588 -15656 14412
rect -14340 14412 -14244 14428
rect -15333 14360 -14611 14361
rect -15333 13640 -15332 14360
rect -14612 13640 -14611 14360
rect -15333 13639 -14611 13640
rect -15752 13572 -15656 13588
rect -14340 13588 -14324 14412
rect -14260 13588 -14244 14412
rect -12928 14412 -12832 14428
rect -13921 14360 -13199 14361
rect -13921 13640 -13920 14360
rect -13200 13640 -13199 14360
rect -13921 13639 -13199 13640
rect -14340 13572 -14244 13588
rect -12928 13588 -12912 14412
rect -12848 13588 -12832 14412
rect -11516 14412 -11420 14428
rect -12509 14360 -11787 14361
rect -12509 13640 -12508 14360
rect -11788 13640 -11787 14360
rect -12509 13639 -11787 13640
rect -12928 13572 -12832 13588
rect -11516 13588 -11500 14412
rect -11436 13588 -11420 14412
rect -10104 14412 -10008 14428
rect -11097 14360 -10375 14361
rect -11097 13640 -11096 14360
rect -10376 13640 -10375 14360
rect -11097 13639 -10375 13640
rect -11516 13572 -11420 13588
rect -10104 13588 -10088 14412
rect -10024 13588 -10008 14412
rect -8692 14412 -8596 14428
rect -9685 14360 -8963 14361
rect -9685 13640 -9684 14360
rect -8964 13640 -8963 14360
rect -9685 13639 -8963 13640
rect -10104 13572 -10008 13588
rect -8692 13588 -8676 14412
rect -8612 13588 -8596 14412
rect -7280 14412 -7184 14428
rect -8273 14360 -7551 14361
rect -8273 13640 -8272 14360
rect -7552 13640 -7551 14360
rect -8273 13639 -7551 13640
rect -8692 13572 -8596 13588
rect -7280 13588 -7264 14412
rect -7200 13588 -7184 14412
rect -5868 14412 -5772 14428
rect -6861 14360 -6139 14361
rect -6861 13640 -6860 14360
rect -6140 13640 -6139 14360
rect -6861 13639 -6139 13640
rect -7280 13572 -7184 13588
rect -5868 13588 -5852 14412
rect -5788 13588 -5772 14412
rect -4456 14412 -4360 14428
rect -5449 14360 -4727 14361
rect -5449 13640 -5448 14360
rect -4728 13640 -4727 14360
rect -5449 13639 -4727 13640
rect -5868 13572 -5772 13588
rect -4456 13588 -4440 14412
rect -4376 13588 -4360 14412
rect -3044 14412 -2948 14428
rect -4037 14360 -3315 14361
rect -4037 13640 -4036 14360
rect -3316 13640 -3315 14360
rect -4037 13639 -3315 13640
rect -4456 13572 -4360 13588
rect -3044 13588 -3028 14412
rect -2964 13588 -2948 14412
rect -1632 14412 -1536 14428
rect -2625 14360 -1903 14361
rect -2625 13640 -2624 14360
rect -1904 13640 -1903 14360
rect -2625 13639 -1903 13640
rect -3044 13572 -2948 13588
rect -1632 13588 -1616 14412
rect -1552 13588 -1536 14412
rect -220 14412 -124 14428
rect -1213 14360 -491 14361
rect -1213 13640 -1212 14360
rect -492 13640 -491 14360
rect -1213 13639 -491 13640
rect -1632 13572 -1536 13588
rect -220 13588 -204 14412
rect -140 13588 -124 14412
rect 1192 14412 1288 14428
rect 199 14360 921 14361
rect 199 13640 200 14360
rect 920 13640 921 14360
rect 199 13639 921 13640
rect -220 13572 -124 13588
rect 1192 13588 1208 14412
rect 1272 13588 1288 14412
rect 2604 14412 2700 14428
rect 1611 14360 2333 14361
rect 1611 13640 1612 14360
rect 2332 13640 2333 14360
rect 1611 13639 2333 13640
rect 1192 13572 1288 13588
rect 2604 13588 2620 14412
rect 2684 13588 2700 14412
rect 4016 14412 4112 14428
rect 3023 14360 3745 14361
rect 3023 13640 3024 14360
rect 3744 13640 3745 14360
rect 3023 13639 3745 13640
rect 2604 13572 2700 13588
rect 4016 13588 4032 14412
rect 4096 13588 4112 14412
rect 5428 14412 5524 14428
rect 4435 14360 5157 14361
rect 4435 13640 4436 14360
rect 5156 13640 5157 14360
rect 4435 13639 5157 13640
rect 4016 13572 4112 13588
rect 5428 13588 5444 14412
rect 5508 13588 5524 14412
rect 6840 14412 6936 14428
rect 5847 14360 6569 14361
rect 5847 13640 5848 14360
rect 6568 13640 6569 14360
rect 5847 13639 6569 13640
rect 5428 13572 5524 13588
rect 6840 13588 6856 14412
rect 6920 13588 6936 14412
rect 8252 14412 8348 14428
rect 7259 14360 7981 14361
rect 7259 13640 7260 14360
rect 7980 13640 7981 14360
rect 7259 13639 7981 13640
rect 6840 13572 6936 13588
rect 8252 13588 8268 14412
rect 8332 13588 8348 14412
rect 9664 14412 9760 14428
rect 8671 14360 9393 14361
rect 8671 13640 8672 14360
rect 9392 13640 9393 14360
rect 8671 13639 9393 13640
rect 8252 13572 8348 13588
rect 9664 13588 9680 14412
rect 9744 13588 9760 14412
rect 11076 14412 11172 14428
rect 10083 14360 10805 14361
rect 10083 13640 10084 14360
rect 10804 13640 10805 14360
rect 10083 13639 10805 13640
rect 9664 13572 9760 13588
rect 11076 13588 11092 14412
rect 11156 13588 11172 14412
rect 12488 14412 12584 14428
rect 11495 14360 12217 14361
rect 11495 13640 11496 14360
rect 12216 13640 12217 14360
rect 11495 13639 12217 13640
rect 11076 13572 11172 13588
rect 12488 13588 12504 14412
rect 12568 13588 12584 14412
rect 13900 14412 13996 14428
rect 12907 14360 13629 14361
rect 12907 13640 12908 14360
rect 13628 13640 13629 14360
rect 12907 13639 13629 13640
rect 12488 13572 12584 13588
rect 13900 13588 13916 14412
rect 13980 13588 13996 14412
rect 15312 14412 15408 14428
rect 14319 14360 15041 14361
rect 14319 13640 14320 14360
rect 15040 13640 15041 14360
rect 14319 13639 15041 13640
rect 13900 13572 13996 13588
rect 15312 13588 15328 14412
rect 15392 13588 15408 14412
rect 16724 14412 16820 14428
rect 15731 14360 16453 14361
rect 15731 13640 15732 14360
rect 16452 13640 16453 14360
rect 15731 13639 16453 13640
rect 15312 13572 15408 13588
rect 16724 13588 16740 14412
rect 16804 13588 16820 14412
rect 18136 14412 18232 14428
rect 17143 14360 17865 14361
rect 17143 13640 17144 14360
rect 17864 13640 17865 14360
rect 17143 13639 17865 13640
rect 16724 13572 16820 13588
rect 18136 13588 18152 14412
rect 18216 13588 18232 14412
rect 19548 14412 19644 14428
rect 18555 14360 19277 14361
rect 18555 13640 18556 14360
rect 19276 13640 19277 14360
rect 18555 13639 19277 13640
rect 18136 13572 18232 13588
rect 19548 13588 19564 14412
rect 19628 13588 19644 14412
rect 20960 14412 21056 14428
rect 19967 14360 20689 14361
rect 19967 13640 19968 14360
rect 20688 13640 20689 14360
rect 19967 13639 20689 13640
rect 19548 13572 19644 13588
rect 20960 13588 20976 14412
rect 21040 13588 21056 14412
rect 22372 14412 22468 14428
rect 21379 14360 22101 14361
rect 21379 13640 21380 14360
rect 22100 13640 22101 14360
rect 21379 13639 22101 13640
rect 20960 13572 21056 13588
rect 22372 13588 22388 14412
rect 22452 13588 22468 14412
rect 23784 14412 23880 14428
rect 22791 14360 23513 14361
rect 22791 13640 22792 14360
rect 23512 13640 23513 14360
rect 22791 13639 23513 13640
rect 22372 13572 22468 13588
rect 23784 13588 23800 14412
rect 23864 13588 23880 14412
rect 23784 13572 23880 13588
rect -22812 13292 -22716 13308
rect -23805 13240 -23083 13241
rect -23805 12520 -23804 13240
rect -23084 12520 -23083 13240
rect -23805 12519 -23083 12520
rect -22812 12468 -22796 13292
rect -22732 12468 -22716 13292
rect -21400 13292 -21304 13308
rect -22393 13240 -21671 13241
rect -22393 12520 -22392 13240
rect -21672 12520 -21671 13240
rect -22393 12519 -21671 12520
rect -22812 12452 -22716 12468
rect -21400 12468 -21384 13292
rect -21320 12468 -21304 13292
rect -19988 13292 -19892 13308
rect -20981 13240 -20259 13241
rect -20981 12520 -20980 13240
rect -20260 12520 -20259 13240
rect -20981 12519 -20259 12520
rect -21400 12452 -21304 12468
rect -19988 12468 -19972 13292
rect -19908 12468 -19892 13292
rect -18576 13292 -18480 13308
rect -19569 13240 -18847 13241
rect -19569 12520 -19568 13240
rect -18848 12520 -18847 13240
rect -19569 12519 -18847 12520
rect -19988 12452 -19892 12468
rect -18576 12468 -18560 13292
rect -18496 12468 -18480 13292
rect -17164 13292 -17068 13308
rect -18157 13240 -17435 13241
rect -18157 12520 -18156 13240
rect -17436 12520 -17435 13240
rect -18157 12519 -17435 12520
rect -18576 12452 -18480 12468
rect -17164 12468 -17148 13292
rect -17084 12468 -17068 13292
rect -15752 13292 -15656 13308
rect -16745 13240 -16023 13241
rect -16745 12520 -16744 13240
rect -16024 12520 -16023 13240
rect -16745 12519 -16023 12520
rect -17164 12452 -17068 12468
rect -15752 12468 -15736 13292
rect -15672 12468 -15656 13292
rect -14340 13292 -14244 13308
rect -15333 13240 -14611 13241
rect -15333 12520 -15332 13240
rect -14612 12520 -14611 13240
rect -15333 12519 -14611 12520
rect -15752 12452 -15656 12468
rect -14340 12468 -14324 13292
rect -14260 12468 -14244 13292
rect -12928 13292 -12832 13308
rect -13921 13240 -13199 13241
rect -13921 12520 -13920 13240
rect -13200 12520 -13199 13240
rect -13921 12519 -13199 12520
rect -14340 12452 -14244 12468
rect -12928 12468 -12912 13292
rect -12848 12468 -12832 13292
rect -11516 13292 -11420 13308
rect -12509 13240 -11787 13241
rect -12509 12520 -12508 13240
rect -11788 12520 -11787 13240
rect -12509 12519 -11787 12520
rect -12928 12452 -12832 12468
rect -11516 12468 -11500 13292
rect -11436 12468 -11420 13292
rect -10104 13292 -10008 13308
rect -11097 13240 -10375 13241
rect -11097 12520 -11096 13240
rect -10376 12520 -10375 13240
rect -11097 12519 -10375 12520
rect -11516 12452 -11420 12468
rect -10104 12468 -10088 13292
rect -10024 12468 -10008 13292
rect -8692 13292 -8596 13308
rect -9685 13240 -8963 13241
rect -9685 12520 -9684 13240
rect -8964 12520 -8963 13240
rect -9685 12519 -8963 12520
rect -10104 12452 -10008 12468
rect -8692 12468 -8676 13292
rect -8612 12468 -8596 13292
rect -7280 13292 -7184 13308
rect -8273 13240 -7551 13241
rect -8273 12520 -8272 13240
rect -7552 12520 -7551 13240
rect -8273 12519 -7551 12520
rect -8692 12452 -8596 12468
rect -7280 12468 -7264 13292
rect -7200 12468 -7184 13292
rect -5868 13292 -5772 13308
rect -6861 13240 -6139 13241
rect -6861 12520 -6860 13240
rect -6140 12520 -6139 13240
rect -6861 12519 -6139 12520
rect -7280 12452 -7184 12468
rect -5868 12468 -5852 13292
rect -5788 12468 -5772 13292
rect -4456 13292 -4360 13308
rect -5449 13240 -4727 13241
rect -5449 12520 -5448 13240
rect -4728 12520 -4727 13240
rect -5449 12519 -4727 12520
rect -5868 12452 -5772 12468
rect -4456 12468 -4440 13292
rect -4376 12468 -4360 13292
rect -3044 13292 -2948 13308
rect -4037 13240 -3315 13241
rect -4037 12520 -4036 13240
rect -3316 12520 -3315 13240
rect -4037 12519 -3315 12520
rect -4456 12452 -4360 12468
rect -3044 12468 -3028 13292
rect -2964 12468 -2948 13292
rect -1632 13292 -1536 13308
rect -2625 13240 -1903 13241
rect -2625 12520 -2624 13240
rect -1904 12520 -1903 13240
rect -2625 12519 -1903 12520
rect -3044 12452 -2948 12468
rect -1632 12468 -1616 13292
rect -1552 12468 -1536 13292
rect -220 13292 -124 13308
rect -1213 13240 -491 13241
rect -1213 12520 -1212 13240
rect -492 12520 -491 13240
rect -1213 12519 -491 12520
rect -1632 12452 -1536 12468
rect -220 12468 -204 13292
rect -140 12468 -124 13292
rect 1192 13292 1288 13308
rect 199 13240 921 13241
rect 199 12520 200 13240
rect 920 12520 921 13240
rect 199 12519 921 12520
rect -220 12452 -124 12468
rect 1192 12468 1208 13292
rect 1272 12468 1288 13292
rect 2604 13292 2700 13308
rect 1611 13240 2333 13241
rect 1611 12520 1612 13240
rect 2332 12520 2333 13240
rect 1611 12519 2333 12520
rect 1192 12452 1288 12468
rect 2604 12468 2620 13292
rect 2684 12468 2700 13292
rect 4016 13292 4112 13308
rect 3023 13240 3745 13241
rect 3023 12520 3024 13240
rect 3744 12520 3745 13240
rect 3023 12519 3745 12520
rect 2604 12452 2700 12468
rect 4016 12468 4032 13292
rect 4096 12468 4112 13292
rect 5428 13292 5524 13308
rect 4435 13240 5157 13241
rect 4435 12520 4436 13240
rect 5156 12520 5157 13240
rect 4435 12519 5157 12520
rect 4016 12452 4112 12468
rect 5428 12468 5444 13292
rect 5508 12468 5524 13292
rect 6840 13292 6936 13308
rect 5847 13240 6569 13241
rect 5847 12520 5848 13240
rect 6568 12520 6569 13240
rect 5847 12519 6569 12520
rect 5428 12452 5524 12468
rect 6840 12468 6856 13292
rect 6920 12468 6936 13292
rect 8252 13292 8348 13308
rect 7259 13240 7981 13241
rect 7259 12520 7260 13240
rect 7980 12520 7981 13240
rect 7259 12519 7981 12520
rect 6840 12452 6936 12468
rect 8252 12468 8268 13292
rect 8332 12468 8348 13292
rect 9664 13292 9760 13308
rect 8671 13240 9393 13241
rect 8671 12520 8672 13240
rect 9392 12520 9393 13240
rect 8671 12519 9393 12520
rect 8252 12452 8348 12468
rect 9664 12468 9680 13292
rect 9744 12468 9760 13292
rect 11076 13292 11172 13308
rect 10083 13240 10805 13241
rect 10083 12520 10084 13240
rect 10804 12520 10805 13240
rect 10083 12519 10805 12520
rect 9664 12452 9760 12468
rect 11076 12468 11092 13292
rect 11156 12468 11172 13292
rect 12488 13292 12584 13308
rect 11495 13240 12217 13241
rect 11495 12520 11496 13240
rect 12216 12520 12217 13240
rect 11495 12519 12217 12520
rect 11076 12452 11172 12468
rect 12488 12468 12504 13292
rect 12568 12468 12584 13292
rect 13900 13292 13996 13308
rect 12907 13240 13629 13241
rect 12907 12520 12908 13240
rect 13628 12520 13629 13240
rect 12907 12519 13629 12520
rect 12488 12452 12584 12468
rect 13900 12468 13916 13292
rect 13980 12468 13996 13292
rect 15312 13292 15408 13308
rect 14319 13240 15041 13241
rect 14319 12520 14320 13240
rect 15040 12520 15041 13240
rect 14319 12519 15041 12520
rect 13900 12452 13996 12468
rect 15312 12468 15328 13292
rect 15392 12468 15408 13292
rect 16724 13292 16820 13308
rect 15731 13240 16453 13241
rect 15731 12520 15732 13240
rect 16452 12520 16453 13240
rect 15731 12519 16453 12520
rect 15312 12452 15408 12468
rect 16724 12468 16740 13292
rect 16804 12468 16820 13292
rect 18136 13292 18232 13308
rect 17143 13240 17865 13241
rect 17143 12520 17144 13240
rect 17864 12520 17865 13240
rect 17143 12519 17865 12520
rect 16724 12452 16820 12468
rect 18136 12468 18152 13292
rect 18216 12468 18232 13292
rect 19548 13292 19644 13308
rect 18555 13240 19277 13241
rect 18555 12520 18556 13240
rect 19276 12520 19277 13240
rect 18555 12519 19277 12520
rect 18136 12452 18232 12468
rect 19548 12468 19564 13292
rect 19628 12468 19644 13292
rect 20960 13292 21056 13308
rect 19967 13240 20689 13241
rect 19967 12520 19968 13240
rect 20688 12520 20689 13240
rect 19967 12519 20689 12520
rect 19548 12452 19644 12468
rect 20960 12468 20976 13292
rect 21040 12468 21056 13292
rect 22372 13292 22468 13308
rect 21379 13240 22101 13241
rect 21379 12520 21380 13240
rect 22100 12520 22101 13240
rect 21379 12519 22101 12520
rect 20960 12452 21056 12468
rect 22372 12468 22388 13292
rect 22452 12468 22468 13292
rect 23784 13292 23880 13308
rect 22791 13240 23513 13241
rect 22791 12520 22792 13240
rect 23512 12520 23513 13240
rect 22791 12519 23513 12520
rect 22372 12452 22468 12468
rect 23784 12468 23800 13292
rect 23864 12468 23880 13292
rect 23784 12452 23880 12468
rect -22812 12172 -22716 12188
rect -23805 12120 -23083 12121
rect -23805 11400 -23804 12120
rect -23084 11400 -23083 12120
rect -23805 11399 -23083 11400
rect -22812 11348 -22796 12172
rect -22732 11348 -22716 12172
rect -21400 12172 -21304 12188
rect -22393 12120 -21671 12121
rect -22393 11400 -22392 12120
rect -21672 11400 -21671 12120
rect -22393 11399 -21671 11400
rect -22812 11332 -22716 11348
rect -21400 11348 -21384 12172
rect -21320 11348 -21304 12172
rect -19988 12172 -19892 12188
rect -20981 12120 -20259 12121
rect -20981 11400 -20980 12120
rect -20260 11400 -20259 12120
rect -20981 11399 -20259 11400
rect -21400 11332 -21304 11348
rect -19988 11348 -19972 12172
rect -19908 11348 -19892 12172
rect -18576 12172 -18480 12188
rect -19569 12120 -18847 12121
rect -19569 11400 -19568 12120
rect -18848 11400 -18847 12120
rect -19569 11399 -18847 11400
rect -19988 11332 -19892 11348
rect -18576 11348 -18560 12172
rect -18496 11348 -18480 12172
rect -17164 12172 -17068 12188
rect -18157 12120 -17435 12121
rect -18157 11400 -18156 12120
rect -17436 11400 -17435 12120
rect -18157 11399 -17435 11400
rect -18576 11332 -18480 11348
rect -17164 11348 -17148 12172
rect -17084 11348 -17068 12172
rect -15752 12172 -15656 12188
rect -16745 12120 -16023 12121
rect -16745 11400 -16744 12120
rect -16024 11400 -16023 12120
rect -16745 11399 -16023 11400
rect -17164 11332 -17068 11348
rect -15752 11348 -15736 12172
rect -15672 11348 -15656 12172
rect -14340 12172 -14244 12188
rect -15333 12120 -14611 12121
rect -15333 11400 -15332 12120
rect -14612 11400 -14611 12120
rect -15333 11399 -14611 11400
rect -15752 11332 -15656 11348
rect -14340 11348 -14324 12172
rect -14260 11348 -14244 12172
rect -12928 12172 -12832 12188
rect -13921 12120 -13199 12121
rect -13921 11400 -13920 12120
rect -13200 11400 -13199 12120
rect -13921 11399 -13199 11400
rect -14340 11332 -14244 11348
rect -12928 11348 -12912 12172
rect -12848 11348 -12832 12172
rect -11516 12172 -11420 12188
rect -12509 12120 -11787 12121
rect -12509 11400 -12508 12120
rect -11788 11400 -11787 12120
rect -12509 11399 -11787 11400
rect -12928 11332 -12832 11348
rect -11516 11348 -11500 12172
rect -11436 11348 -11420 12172
rect -10104 12172 -10008 12188
rect -11097 12120 -10375 12121
rect -11097 11400 -11096 12120
rect -10376 11400 -10375 12120
rect -11097 11399 -10375 11400
rect -11516 11332 -11420 11348
rect -10104 11348 -10088 12172
rect -10024 11348 -10008 12172
rect -8692 12172 -8596 12188
rect -9685 12120 -8963 12121
rect -9685 11400 -9684 12120
rect -8964 11400 -8963 12120
rect -9685 11399 -8963 11400
rect -10104 11332 -10008 11348
rect -8692 11348 -8676 12172
rect -8612 11348 -8596 12172
rect -7280 12172 -7184 12188
rect -8273 12120 -7551 12121
rect -8273 11400 -8272 12120
rect -7552 11400 -7551 12120
rect -8273 11399 -7551 11400
rect -8692 11332 -8596 11348
rect -7280 11348 -7264 12172
rect -7200 11348 -7184 12172
rect -5868 12172 -5772 12188
rect -6861 12120 -6139 12121
rect -6861 11400 -6860 12120
rect -6140 11400 -6139 12120
rect -6861 11399 -6139 11400
rect -7280 11332 -7184 11348
rect -5868 11348 -5852 12172
rect -5788 11348 -5772 12172
rect -4456 12172 -4360 12188
rect -5449 12120 -4727 12121
rect -5449 11400 -5448 12120
rect -4728 11400 -4727 12120
rect -5449 11399 -4727 11400
rect -5868 11332 -5772 11348
rect -4456 11348 -4440 12172
rect -4376 11348 -4360 12172
rect -3044 12172 -2948 12188
rect -4037 12120 -3315 12121
rect -4037 11400 -4036 12120
rect -3316 11400 -3315 12120
rect -4037 11399 -3315 11400
rect -4456 11332 -4360 11348
rect -3044 11348 -3028 12172
rect -2964 11348 -2948 12172
rect -1632 12172 -1536 12188
rect -2625 12120 -1903 12121
rect -2625 11400 -2624 12120
rect -1904 11400 -1903 12120
rect -2625 11399 -1903 11400
rect -3044 11332 -2948 11348
rect -1632 11348 -1616 12172
rect -1552 11348 -1536 12172
rect -220 12172 -124 12188
rect -1213 12120 -491 12121
rect -1213 11400 -1212 12120
rect -492 11400 -491 12120
rect -1213 11399 -491 11400
rect -1632 11332 -1536 11348
rect -220 11348 -204 12172
rect -140 11348 -124 12172
rect 1192 12172 1288 12188
rect 199 12120 921 12121
rect 199 11400 200 12120
rect 920 11400 921 12120
rect 199 11399 921 11400
rect -220 11332 -124 11348
rect 1192 11348 1208 12172
rect 1272 11348 1288 12172
rect 2604 12172 2700 12188
rect 1611 12120 2333 12121
rect 1611 11400 1612 12120
rect 2332 11400 2333 12120
rect 1611 11399 2333 11400
rect 1192 11332 1288 11348
rect 2604 11348 2620 12172
rect 2684 11348 2700 12172
rect 4016 12172 4112 12188
rect 3023 12120 3745 12121
rect 3023 11400 3024 12120
rect 3744 11400 3745 12120
rect 3023 11399 3745 11400
rect 2604 11332 2700 11348
rect 4016 11348 4032 12172
rect 4096 11348 4112 12172
rect 5428 12172 5524 12188
rect 4435 12120 5157 12121
rect 4435 11400 4436 12120
rect 5156 11400 5157 12120
rect 4435 11399 5157 11400
rect 4016 11332 4112 11348
rect 5428 11348 5444 12172
rect 5508 11348 5524 12172
rect 6840 12172 6936 12188
rect 5847 12120 6569 12121
rect 5847 11400 5848 12120
rect 6568 11400 6569 12120
rect 5847 11399 6569 11400
rect 5428 11332 5524 11348
rect 6840 11348 6856 12172
rect 6920 11348 6936 12172
rect 8252 12172 8348 12188
rect 7259 12120 7981 12121
rect 7259 11400 7260 12120
rect 7980 11400 7981 12120
rect 7259 11399 7981 11400
rect 6840 11332 6936 11348
rect 8252 11348 8268 12172
rect 8332 11348 8348 12172
rect 9664 12172 9760 12188
rect 8671 12120 9393 12121
rect 8671 11400 8672 12120
rect 9392 11400 9393 12120
rect 8671 11399 9393 11400
rect 8252 11332 8348 11348
rect 9664 11348 9680 12172
rect 9744 11348 9760 12172
rect 11076 12172 11172 12188
rect 10083 12120 10805 12121
rect 10083 11400 10084 12120
rect 10804 11400 10805 12120
rect 10083 11399 10805 11400
rect 9664 11332 9760 11348
rect 11076 11348 11092 12172
rect 11156 11348 11172 12172
rect 12488 12172 12584 12188
rect 11495 12120 12217 12121
rect 11495 11400 11496 12120
rect 12216 11400 12217 12120
rect 11495 11399 12217 11400
rect 11076 11332 11172 11348
rect 12488 11348 12504 12172
rect 12568 11348 12584 12172
rect 13900 12172 13996 12188
rect 12907 12120 13629 12121
rect 12907 11400 12908 12120
rect 13628 11400 13629 12120
rect 12907 11399 13629 11400
rect 12488 11332 12584 11348
rect 13900 11348 13916 12172
rect 13980 11348 13996 12172
rect 15312 12172 15408 12188
rect 14319 12120 15041 12121
rect 14319 11400 14320 12120
rect 15040 11400 15041 12120
rect 14319 11399 15041 11400
rect 13900 11332 13996 11348
rect 15312 11348 15328 12172
rect 15392 11348 15408 12172
rect 16724 12172 16820 12188
rect 15731 12120 16453 12121
rect 15731 11400 15732 12120
rect 16452 11400 16453 12120
rect 15731 11399 16453 11400
rect 15312 11332 15408 11348
rect 16724 11348 16740 12172
rect 16804 11348 16820 12172
rect 18136 12172 18232 12188
rect 17143 12120 17865 12121
rect 17143 11400 17144 12120
rect 17864 11400 17865 12120
rect 17143 11399 17865 11400
rect 16724 11332 16820 11348
rect 18136 11348 18152 12172
rect 18216 11348 18232 12172
rect 19548 12172 19644 12188
rect 18555 12120 19277 12121
rect 18555 11400 18556 12120
rect 19276 11400 19277 12120
rect 18555 11399 19277 11400
rect 18136 11332 18232 11348
rect 19548 11348 19564 12172
rect 19628 11348 19644 12172
rect 20960 12172 21056 12188
rect 19967 12120 20689 12121
rect 19967 11400 19968 12120
rect 20688 11400 20689 12120
rect 19967 11399 20689 11400
rect 19548 11332 19644 11348
rect 20960 11348 20976 12172
rect 21040 11348 21056 12172
rect 22372 12172 22468 12188
rect 21379 12120 22101 12121
rect 21379 11400 21380 12120
rect 22100 11400 22101 12120
rect 21379 11399 22101 11400
rect 20960 11332 21056 11348
rect 22372 11348 22388 12172
rect 22452 11348 22468 12172
rect 23784 12172 23880 12188
rect 22791 12120 23513 12121
rect 22791 11400 22792 12120
rect 23512 11400 23513 12120
rect 22791 11399 23513 11400
rect 22372 11332 22468 11348
rect 23784 11348 23800 12172
rect 23864 11348 23880 12172
rect 23784 11332 23880 11348
rect -22812 11052 -22716 11068
rect -23805 11000 -23083 11001
rect -23805 10280 -23804 11000
rect -23084 10280 -23083 11000
rect -23805 10279 -23083 10280
rect -22812 10228 -22796 11052
rect -22732 10228 -22716 11052
rect -21400 11052 -21304 11068
rect -22393 11000 -21671 11001
rect -22393 10280 -22392 11000
rect -21672 10280 -21671 11000
rect -22393 10279 -21671 10280
rect -22812 10212 -22716 10228
rect -21400 10228 -21384 11052
rect -21320 10228 -21304 11052
rect -19988 11052 -19892 11068
rect -20981 11000 -20259 11001
rect -20981 10280 -20980 11000
rect -20260 10280 -20259 11000
rect -20981 10279 -20259 10280
rect -21400 10212 -21304 10228
rect -19988 10228 -19972 11052
rect -19908 10228 -19892 11052
rect -18576 11052 -18480 11068
rect -19569 11000 -18847 11001
rect -19569 10280 -19568 11000
rect -18848 10280 -18847 11000
rect -19569 10279 -18847 10280
rect -19988 10212 -19892 10228
rect -18576 10228 -18560 11052
rect -18496 10228 -18480 11052
rect -17164 11052 -17068 11068
rect -18157 11000 -17435 11001
rect -18157 10280 -18156 11000
rect -17436 10280 -17435 11000
rect -18157 10279 -17435 10280
rect -18576 10212 -18480 10228
rect -17164 10228 -17148 11052
rect -17084 10228 -17068 11052
rect -15752 11052 -15656 11068
rect -16745 11000 -16023 11001
rect -16745 10280 -16744 11000
rect -16024 10280 -16023 11000
rect -16745 10279 -16023 10280
rect -17164 10212 -17068 10228
rect -15752 10228 -15736 11052
rect -15672 10228 -15656 11052
rect -14340 11052 -14244 11068
rect -15333 11000 -14611 11001
rect -15333 10280 -15332 11000
rect -14612 10280 -14611 11000
rect -15333 10279 -14611 10280
rect -15752 10212 -15656 10228
rect -14340 10228 -14324 11052
rect -14260 10228 -14244 11052
rect -12928 11052 -12832 11068
rect -13921 11000 -13199 11001
rect -13921 10280 -13920 11000
rect -13200 10280 -13199 11000
rect -13921 10279 -13199 10280
rect -14340 10212 -14244 10228
rect -12928 10228 -12912 11052
rect -12848 10228 -12832 11052
rect -11516 11052 -11420 11068
rect -12509 11000 -11787 11001
rect -12509 10280 -12508 11000
rect -11788 10280 -11787 11000
rect -12509 10279 -11787 10280
rect -12928 10212 -12832 10228
rect -11516 10228 -11500 11052
rect -11436 10228 -11420 11052
rect -10104 11052 -10008 11068
rect -11097 11000 -10375 11001
rect -11097 10280 -11096 11000
rect -10376 10280 -10375 11000
rect -11097 10279 -10375 10280
rect -11516 10212 -11420 10228
rect -10104 10228 -10088 11052
rect -10024 10228 -10008 11052
rect -8692 11052 -8596 11068
rect -9685 11000 -8963 11001
rect -9685 10280 -9684 11000
rect -8964 10280 -8963 11000
rect -9685 10279 -8963 10280
rect -10104 10212 -10008 10228
rect -8692 10228 -8676 11052
rect -8612 10228 -8596 11052
rect -7280 11052 -7184 11068
rect -8273 11000 -7551 11001
rect -8273 10280 -8272 11000
rect -7552 10280 -7551 11000
rect -8273 10279 -7551 10280
rect -8692 10212 -8596 10228
rect -7280 10228 -7264 11052
rect -7200 10228 -7184 11052
rect -5868 11052 -5772 11068
rect -6861 11000 -6139 11001
rect -6861 10280 -6860 11000
rect -6140 10280 -6139 11000
rect -6861 10279 -6139 10280
rect -7280 10212 -7184 10228
rect -5868 10228 -5852 11052
rect -5788 10228 -5772 11052
rect -4456 11052 -4360 11068
rect -5449 11000 -4727 11001
rect -5449 10280 -5448 11000
rect -4728 10280 -4727 11000
rect -5449 10279 -4727 10280
rect -5868 10212 -5772 10228
rect -4456 10228 -4440 11052
rect -4376 10228 -4360 11052
rect -3044 11052 -2948 11068
rect -4037 11000 -3315 11001
rect -4037 10280 -4036 11000
rect -3316 10280 -3315 11000
rect -4037 10279 -3315 10280
rect -4456 10212 -4360 10228
rect -3044 10228 -3028 11052
rect -2964 10228 -2948 11052
rect -1632 11052 -1536 11068
rect -2625 11000 -1903 11001
rect -2625 10280 -2624 11000
rect -1904 10280 -1903 11000
rect -2625 10279 -1903 10280
rect -3044 10212 -2948 10228
rect -1632 10228 -1616 11052
rect -1552 10228 -1536 11052
rect -220 11052 -124 11068
rect -1213 11000 -491 11001
rect -1213 10280 -1212 11000
rect -492 10280 -491 11000
rect -1213 10279 -491 10280
rect -1632 10212 -1536 10228
rect -220 10228 -204 11052
rect -140 10228 -124 11052
rect 1192 11052 1288 11068
rect 199 11000 921 11001
rect 199 10280 200 11000
rect 920 10280 921 11000
rect 199 10279 921 10280
rect -220 10212 -124 10228
rect 1192 10228 1208 11052
rect 1272 10228 1288 11052
rect 2604 11052 2700 11068
rect 1611 11000 2333 11001
rect 1611 10280 1612 11000
rect 2332 10280 2333 11000
rect 1611 10279 2333 10280
rect 1192 10212 1288 10228
rect 2604 10228 2620 11052
rect 2684 10228 2700 11052
rect 4016 11052 4112 11068
rect 3023 11000 3745 11001
rect 3023 10280 3024 11000
rect 3744 10280 3745 11000
rect 3023 10279 3745 10280
rect 2604 10212 2700 10228
rect 4016 10228 4032 11052
rect 4096 10228 4112 11052
rect 5428 11052 5524 11068
rect 4435 11000 5157 11001
rect 4435 10280 4436 11000
rect 5156 10280 5157 11000
rect 4435 10279 5157 10280
rect 4016 10212 4112 10228
rect 5428 10228 5444 11052
rect 5508 10228 5524 11052
rect 6840 11052 6936 11068
rect 5847 11000 6569 11001
rect 5847 10280 5848 11000
rect 6568 10280 6569 11000
rect 5847 10279 6569 10280
rect 5428 10212 5524 10228
rect 6840 10228 6856 11052
rect 6920 10228 6936 11052
rect 8252 11052 8348 11068
rect 7259 11000 7981 11001
rect 7259 10280 7260 11000
rect 7980 10280 7981 11000
rect 7259 10279 7981 10280
rect 6840 10212 6936 10228
rect 8252 10228 8268 11052
rect 8332 10228 8348 11052
rect 9664 11052 9760 11068
rect 8671 11000 9393 11001
rect 8671 10280 8672 11000
rect 9392 10280 9393 11000
rect 8671 10279 9393 10280
rect 8252 10212 8348 10228
rect 9664 10228 9680 11052
rect 9744 10228 9760 11052
rect 11076 11052 11172 11068
rect 10083 11000 10805 11001
rect 10083 10280 10084 11000
rect 10804 10280 10805 11000
rect 10083 10279 10805 10280
rect 9664 10212 9760 10228
rect 11076 10228 11092 11052
rect 11156 10228 11172 11052
rect 12488 11052 12584 11068
rect 11495 11000 12217 11001
rect 11495 10280 11496 11000
rect 12216 10280 12217 11000
rect 11495 10279 12217 10280
rect 11076 10212 11172 10228
rect 12488 10228 12504 11052
rect 12568 10228 12584 11052
rect 13900 11052 13996 11068
rect 12907 11000 13629 11001
rect 12907 10280 12908 11000
rect 13628 10280 13629 11000
rect 12907 10279 13629 10280
rect 12488 10212 12584 10228
rect 13900 10228 13916 11052
rect 13980 10228 13996 11052
rect 15312 11052 15408 11068
rect 14319 11000 15041 11001
rect 14319 10280 14320 11000
rect 15040 10280 15041 11000
rect 14319 10279 15041 10280
rect 13900 10212 13996 10228
rect 15312 10228 15328 11052
rect 15392 10228 15408 11052
rect 16724 11052 16820 11068
rect 15731 11000 16453 11001
rect 15731 10280 15732 11000
rect 16452 10280 16453 11000
rect 15731 10279 16453 10280
rect 15312 10212 15408 10228
rect 16724 10228 16740 11052
rect 16804 10228 16820 11052
rect 18136 11052 18232 11068
rect 17143 11000 17865 11001
rect 17143 10280 17144 11000
rect 17864 10280 17865 11000
rect 17143 10279 17865 10280
rect 16724 10212 16820 10228
rect 18136 10228 18152 11052
rect 18216 10228 18232 11052
rect 19548 11052 19644 11068
rect 18555 11000 19277 11001
rect 18555 10280 18556 11000
rect 19276 10280 19277 11000
rect 18555 10279 19277 10280
rect 18136 10212 18232 10228
rect 19548 10228 19564 11052
rect 19628 10228 19644 11052
rect 20960 11052 21056 11068
rect 19967 11000 20689 11001
rect 19967 10280 19968 11000
rect 20688 10280 20689 11000
rect 19967 10279 20689 10280
rect 19548 10212 19644 10228
rect 20960 10228 20976 11052
rect 21040 10228 21056 11052
rect 22372 11052 22468 11068
rect 21379 11000 22101 11001
rect 21379 10280 21380 11000
rect 22100 10280 22101 11000
rect 21379 10279 22101 10280
rect 20960 10212 21056 10228
rect 22372 10228 22388 11052
rect 22452 10228 22468 11052
rect 23784 11052 23880 11068
rect 22791 11000 23513 11001
rect 22791 10280 22792 11000
rect 23512 10280 23513 11000
rect 22791 10279 23513 10280
rect 22372 10212 22468 10228
rect 23784 10228 23800 11052
rect 23864 10228 23880 11052
rect 23784 10212 23880 10228
rect -22812 9932 -22716 9948
rect -23805 9880 -23083 9881
rect -23805 9160 -23804 9880
rect -23084 9160 -23083 9880
rect -23805 9159 -23083 9160
rect -22812 9108 -22796 9932
rect -22732 9108 -22716 9932
rect -21400 9932 -21304 9948
rect -22393 9880 -21671 9881
rect -22393 9160 -22392 9880
rect -21672 9160 -21671 9880
rect -22393 9159 -21671 9160
rect -22812 9092 -22716 9108
rect -21400 9108 -21384 9932
rect -21320 9108 -21304 9932
rect -19988 9932 -19892 9948
rect -20981 9880 -20259 9881
rect -20981 9160 -20980 9880
rect -20260 9160 -20259 9880
rect -20981 9159 -20259 9160
rect -21400 9092 -21304 9108
rect -19988 9108 -19972 9932
rect -19908 9108 -19892 9932
rect -18576 9932 -18480 9948
rect -19569 9880 -18847 9881
rect -19569 9160 -19568 9880
rect -18848 9160 -18847 9880
rect -19569 9159 -18847 9160
rect -19988 9092 -19892 9108
rect -18576 9108 -18560 9932
rect -18496 9108 -18480 9932
rect -17164 9932 -17068 9948
rect -18157 9880 -17435 9881
rect -18157 9160 -18156 9880
rect -17436 9160 -17435 9880
rect -18157 9159 -17435 9160
rect -18576 9092 -18480 9108
rect -17164 9108 -17148 9932
rect -17084 9108 -17068 9932
rect -15752 9932 -15656 9948
rect -16745 9880 -16023 9881
rect -16745 9160 -16744 9880
rect -16024 9160 -16023 9880
rect -16745 9159 -16023 9160
rect -17164 9092 -17068 9108
rect -15752 9108 -15736 9932
rect -15672 9108 -15656 9932
rect -14340 9932 -14244 9948
rect -15333 9880 -14611 9881
rect -15333 9160 -15332 9880
rect -14612 9160 -14611 9880
rect -15333 9159 -14611 9160
rect -15752 9092 -15656 9108
rect -14340 9108 -14324 9932
rect -14260 9108 -14244 9932
rect -12928 9932 -12832 9948
rect -13921 9880 -13199 9881
rect -13921 9160 -13920 9880
rect -13200 9160 -13199 9880
rect -13921 9159 -13199 9160
rect -14340 9092 -14244 9108
rect -12928 9108 -12912 9932
rect -12848 9108 -12832 9932
rect -11516 9932 -11420 9948
rect -12509 9880 -11787 9881
rect -12509 9160 -12508 9880
rect -11788 9160 -11787 9880
rect -12509 9159 -11787 9160
rect -12928 9092 -12832 9108
rect -11516 9108 -11500 9932
rect -11436 9108 -11420 9932
rect -10104 9932 -10008 9948
rect -11097 9880 -10375 9881
rect -11097 9160 -11096 9880
rect -10376 9160 -10375 9880
rect -11097 9159 -10375 9160
rect -11516 9092 -11420 9108
rect -10104 9108 -10088 9932
rect -10024 9108 -10008 9932
rect -8692 9932 -8596 9948
rect -9685 9880 -8963 9881
rect -9685 9160 -9684 9880
rect -8964 9160 -8963 9880
rect -9685 9159 -8963 9160
rect -10104 9092 -10008 9108
rect -8692 9108 -8676 9932
rect -8612 9108 -8596 9932
rect -7280 9932 -7184 9948
rect -8273 9880 -7551 9881
rect -8273 9160 -8272 9880
rect -7552 9160 -7551 9880
rect -8273 9159 -7551 9160
rect -8692 9092 -8596 9108
rect -7280 9108 -7264 9932
rect -7200 9108 -7184 9932
rect -5868 9932 -5772 9948
rect -6861 9880 -6139 9881
rect -6861 9160 -6860 9880
rect -6140 9160 -6139 9880
rect -6861 9159 -6139 9160
rect -7280 9092 -7184 9108
rect -5868 9108 -5852 9932
rect -5788 9108 -5772 9932
rect -4456 9932 -4360 9948
rect -5449 9880 -4727 9881
rect -5449 9160 -5448 9880
rect -4728 9160 -4727 9880
rect -5449 9159 -4727 9160
rect -5868 9092 -5772 9108
rect -4456 9108 -4440 9932
rect -4376 9108 -4360 9932
rect -3044 9932 -2948 9948
rect -4037 9880 -3315 9881
rect -4037 9160 -4036 9880
rect -3316 9160 -3315 9880
rect -4037 9159 -3315 9160
rect -4456 9092 -4360 9108
rect -3044 9108 -3028 9932
rect -2964 9108 -2948 9932
rect -1632 9932 -1536 9948
rect -2625 9880 -1903 9881
rect -2625 9160 -2624 9880
rect -1904 9160 -1903 9880
rect -2625 9159 -1903 9160
rect -3044 9092 -2948 9108
rect -1632 9108 -1616 9932
rect -1552 9108 -1536 9932
rect -220 9932 -124 9948
rect -1213 9880 -491 9881
rect -1213 9160 -1212 9880
rect -492 9160 -491 9880
rect -1213 9159 -491 9160
rect -1632 9092 -1536 9108
rect -220 9108 -204 9932
rect -140 9108 -124 9932
rect 1192 9932 1288 9948
rect 199 9880 921 9881
rect 199 9160 200 9880
rect 920 9160 921 9880
rect 199 9159 921 9160
rect -220 9092 -124 9108
rect 1192 9108 1208 9932
rect 1272 9108 1288 9932
rect 2604 9932 2700 9948
rect 1611 9880 2333 9881
rect 1611 9160 1612 9880
rect 2332 9160 2333 9880
rect 1611 9159 2333 9160
rect 1192 9092 1288 9108
rect 2604 9108 2620 9932
rect 2684 9108 2700 9932
rect 4016 9932 4112 9948
rect 3023 9880 3745 9881
rect 3023 9160 3024 9880
rect 3744 9160 3745 9880
rect 3023 9159 3745 9160
rect 2604 9092 2700 9108
rect 4016 9108 4032 9932
rect 4096 9108 4112 9932
rect 5428 9932 5524 9948
rect 4435 9880 5157 9881
rect 4435 9160 4436 9880
rect 5156 9160 5157 9880
rect 4435 9159 5157 9160
rect 4016 9092 4112 9108
rect 5428 9108 5444 9932
rect 5508 9108 5524 9932
rect 6840 9932 6936 9948
rect 5847 9880 6569 9881
rect 5847 9160 5848 9880
rect 6568 9160 6569 9880
rect 5847 9159 6569 9160
rect 5428 9092 5524 9108
rect 6840 9108 6856 9932
rect 6920 9108 6936 9932
rect 8252 9932 8348 9948
rect 7259 9880 7981 9881
rect 7259 9160 7260 9880
rect 7980 9160 7981 9880
rect 7259 9159 7981 9160
rect 6840 9092 6936 9108
rect 8252 9108 8268 9932
rect 8332 9108 8348 9932
rect 9664 9932 9760 9948
rect 8671 9880 9393 9881
rect 8671 9160 8672 9880
rect 9392 9160 9393 9880
rect 8671 9159 9393 9160
rect 8252 9092 8348 9108
rect 9664 9108 9680 9932
rect 9744 9108 9760 9932
rect 11076 9932 11172 9948
rect 10083 9880 10805 9881
rect 10083 9160 10084 9880
rect 10804 9160 10805 9880
rect 10083 9159 10805 9160
rect 9664 9092 9760 9108
rect 11076 9108 11092 9932
rect 11156 9108 11172 9932
rect 12488 9932 12584 9948
rect 11495 9880 12217 9881
rect 11495 9160 11496 9880
rect 12216 9160 12217 9880
rect 11495 9159 12217 9160
rect 11076 9092 11172 9108
rect 12488 9108 12504 9932
rect 12568 9108 12584 9932
rect 13900 9932 13996 9948
rect 12907 9880 13629 9881
rect 12907 9160 12908 9880
rect 13628 9160 13629 9880
rect 12907 9159 13629 9160
rect 12488 9092 12584 9108
rect 13900 9108 13916 9932
rect 13980 9108 13996 9932
rect 15312 9932 15408 9948
rect 14319 9880 15041 9881
rect 14319 9160 14320 9880
rect 15040 9160 15041 9880
rect 14319 9159 15041 9160
rect 13900 9092 13996 9108
rect 15312 9108 15328 9932
rect 15392 9108 15408 9932
rect 16724 9932 16820 9948
rect 15731 9880 16453 9881
rect 15731 9160 15732 9880
rect 16452 9160 16453 9880
rect 15731 9159 16453 9160
rect 15312 9092 15408 9108
rect 16724 9108 16740 9932
rect 16804 9108 16820 9932
rect 18136 9932 18232 9948
rect 17143 9880 17865 9881
rect 17143 9160 17144 9880
rect 17864 9160 17865 9880
rect 17143 9159 17865 9160
rect 16724 9092 16820 9108
rect 18136 9108 18152 9932
rect 18216 9108 18232 9932
rect 19548 9932 19644 9948
rect 18555 9880 19277 9881
rect 18555 9160 18556 9880
rect 19276 9160 19277 9880
rect 18555 9159 19277 9160
rect 18136 9092 18232 9108
rect 19548 9108 19564 9932
rect 19628 9108 19644 9932
rect 20960 9932 21056 9948
rect 19967 9880 20689 9881
rect 19967 9160 19968 9880
rect 20688 9160 20689 9880
rect 19967 9159 20689 9160
rect 19548 9092 19644 9108
rect 20960 9108 20976 9932
rect 21040 9108 21056 9932
rect 22372 9932 22468 9948
rect 21379 9880 22101 9881
rect 21379 9160 21380 9880
rect 22100 9160 22101 9880
rect 21379 9159 22101 9160
rect 20960 9092 21056 9108
rect 22372 9108 22388 9932
rect 22452 9108 22468 9932
rect 23784 9932 23880 9948
rect 22791 9880 23513 9881
rect 22791 9160 22792 9880
rect 23512 9160 23513 9880
rect 22791 9159 23513 9160
rect 22372 9092 22468 9108
rect 23784 9108 23800 9932
rect 23864 9108 23880 9932
rect 23784 9092 23880 9108
rect -22812 8812 -22716 8828
rect -23805 8760 -23083 8761
rect -23805 8040 -23804 8760
rect -23084 8040 -23083 8760
rect -23805 8039 -23083 8040
rect -22812 7988 -22796 8812
rect -22732 7988 -22716 8812
rect -21400 8812 -21304 8828
rect -22393 8760 -21671 8761
rect -22393 8040 -22392 8760
rect -21672 8040 -21671 8760
rect -22393 8039 -21671 8040
rect -22812 7972 -22716 7988
rect -21400 7988 -21384 8812
rect -21320 7988 -21304 8812
rect -19988 8812 -19892 8828
rect -20981 8760 -20259 8761
rect -20981 8040 -20980 8760
rect -20260 8040 -20259 8760
rect -20981 8039 -20259 8040
rect -21400 7972 -21304 7988
rect -19988 7988 -19972 8812
rect -19908 7988 -19892 8812
rect -18576 8812 -18480 8828
rect -19569 8760 -18847 8761
rect -19569 8040 -19568 8760
rect -18848 8040 -18847 8760
rect -19569 8039 -18847 8040
rect -19988 7972 -19892 7988
rect -18576 7988 -18560 8812
rect -18496 7988 -18480 8812
rect -17164 8812 -17068 8828
rect -18157 8760 -17435 8761
rect -18157 8040 -18156 8760
rect -17436 8040 -17435 8760
rect -18157 8039 -17435 8040
rect -18576 7972 -18480 7988
rect -17164 7988 -17148 8812
rect -17084 7988 -17068 8812
rect -15752 8812 -15656 8828
rect -16745 8760 -16023 8761
rect -16745 8040 -16744 8760
rect -16024 8040 -16023 8760
rect -16745 8039 -16023 8040
rect -17164 7972 -17068 7988
rect -15752 7988 -15736 8812
rect -15672 7988 -15656 8812
rect -14340 8812 -14244 8828
rect -15333 8760 -14611 8761
rect -15333 8040 -15332 8760
rect -14612 8040 -14611 8760
rect -15333 8039 -14611 8040
rect -15752 7972 -15656 7988
rect -14340 7988 -14324 8812
rect -14260 7988 -14244 8812
rect -12928 8812 -12832 8828
rect -13921 8760 -13199 8761
rect -13921 8040 -13920 8760
rect -13200 8040 -13199 8760
rect -13921 8039 -13199 8040
rect -14340 7972 -14244 7988
rect -12928 7988 -12912 8812
rect -12848 7988 -12832 8812
rect -11516 8812 -11420 8828
rect -12509 8760 -11787 8761
rect -12509 8040 -12508 8760
rect -11788 8040 -11787 8760
rect -12509 8039 -11787 8040
rect -12928 7972 -12832 7988
rect -11516 7988 -11500 8812
rect -11436 7988 -11420 8812
rect -10104 8812 -10008 8828
rect -11097 8760 -10375 8761
rect -11097 8040 -11096 8760
rect -10376 8040 -10375 8760
rect -11097 8039 -10375 8040
rect -11516 7972 -11420 7988
rect -10104 7988 -10088 8812
rect -10024 7988 -10008 8812
rect -8692 8812 -8596 8828
rect -9685 8760 -8963 8761
rect -9685 8040 -9684 8760
rect -8964 8040 -8963 8760
rect -9685 8039 -8963 8040
rect -10104 7972 -10008 7988
rect -8692 7988 -8676 8812
rect -8612 7988 -8596 8812
rect -7280 8812 -7184 8828
rect -8273 8760 -7551 8761
rect -8273 8040 -8272 8760
rect -7552 8040 -7551 8760
rect -8273 8039 -7551 8040
rect -8692 7972 -8596 7988
rect -7280 7988 -7264 8812
rect -7200 7988 -7184 8812
rect -5868 8812 -5772 8828
rect -6861 8760 -6139 8761
rect -6861 8040 -6860 8760
rect -6140 8040 -6139 8760
rect -6861 8039 -6139 8040
rect -7280 7972 -7184 7988
rect -5868 7988 -5852 8812
rect -5788 7988 -5772 8812
rect -4456 8812 -4360 8828
rect -5449 8760 -4727 8761
rect -5449 8040 -5448 8760
rect -4728 8040 -4727 8760
rect -5449 8039 -4727 8040
rect -5868 7972 -5772 7988
rect -4456 7988 -4440 8812
rect -4376 7988 -4360 8812
rect -3044 8812 -2948 8828
rect -4037 8760 -3315 8761
rect -4037 8040 -4036 8760
rect -3316 8040 -3315 8760
rect -4037 8039 -3315 8040
rect -4456 7972 -4360 7988
rect -3044 7988 -3028 8812
rect -2964 7988 -2948 8812
rect -1632 8812 -1536 8828
rect -2625 8760 -1903 8761
rect -2625 8040 -2624 8760
rect -1904 8040 -1903 8760
rect -2625 8039 -1903 8040
rect -3044 7972 -2948 7988
rect -1632 7988 -1616 8812
rect -1552 7988 -1536 8812
rect -220 8812 -124 8828
rect -1213 8760 -491 8761
rect -1213 8040 -1212 8760
rect -492 8040 -491 8760
rect -1213 8039 -491 8040
rect -1632 7972 -1536 7988
rect -220 7988 -204 8812
rect -140 7988 -124 8812
rect 1192 8812 1288 8828
rect 199 8760 921 8761
rect 199 8040 200 8760
rect 920 8040 921 8760
rect 199 8039 921 8040
rect -220 7972 -124 7988
rect 1192 7988 1208 8812
rect 1272 7988 1288 8812
rect 2604 8812 2700 8828
rect 1611 8760 2333 8761
rect 1611 8040 1612 8760
rect 2332 8040 2333 8760
rect 1611 8039 2333 8040
rect 1192 7972 1288 7988
rect 2604 7988 2620 8812
rect 2684 7988 2700 8812
rect 4016 8812 4112 8828
rect 3023 8760 3745 8761
rect 3023 8040 3024 8760
rect 3744 8040 3745 8760
rect 3023 8039 3745 8040
rect 2604 7972 2700 7988
rect 4016 7988 4032 8812
rect 4096 7988 4112 8812
rect 5428 8812 5524 8828
rect 4435 8760 5157 8761
rect 4435 8040 4436 8760
rect 5156 8040 5157 8760
rect 4435 8039 5157 8040
rect 4016 7972 4112 7988
rect 5428 7988 5444 8812
rect 5508 7988 5524 8812
rect 6840 8812 6936 8828
rect 5847 8760 6569 8761
rect 5847 8040 5848 8760
rect 6568 8040 6569 8760
rect 5847 8039 6569 8040
rect 5428 7972 5524 7988
rect 6840 7988 6856 8812
rect 6920 7988 6936 8812
rect 8252 8812 8348 8828
rect 7259 8760 7981 8761
rect 7259 8040 7260 8760
rect 7980 8040 7981 8760
rect 7259 8039 7981 8040
rect 6840 7972 6936 7988
rect 8252 7988 8268 8812
rect 8332 7988 8348 8812
rect 9664 8812 9760 8828
rect 8671 8760 9393 8761
rect 8671 8040 8672 8760
rect 9392 8040 9393 8760
rect 8671 8039 9393 8040
rect 8252 7972 8348 7988
rect 9664 7988 9680 8812
rect 9744 7988 9760 8812
rect 11076 8812 11172 8828
rect 10083 8760 10805 8761
rect 10083 8040 10084 8760
rect 10804 8040 10805 8760
rect 10083 8039 10805 8040
rect 9664 7972 9760 7988
rect 11076 7988 11092 8812
rect 11156 7988 11172 8812
rect 12488 8812 12584 8828
rect 11495 8760 12217 8761
rect 11495 8040 11496 8760
rect 12216 8040 12217 8760
rect 11495 8039 12217 8040
rect 11076 7972 11172 7988
rect 12488 7988 12504 8812
rect 12568 7988 12584 8812
rect 13900 8812 13996 8828
rect 12907 8760 13629 8761
rect 12907 8040 12908 8760
rect 13628 8040 13629 8760
rect 12907 8039 13629 8040
rect 12488 7972 12584 7988
rect 13900 7988 13916 8812
rect 13980 7988 13996 8812
rect 15312 8812 15408 8828
rect 14319 8760 15041 8761
rect 14319 8040 14320 8760
rect 15040 8040 15041 8760
rect 14319 8039 15041 8040
rect 13900 7972 13996 7988
rect 15312 7988 15328 8812
rect 15392 7988 15408 8812
rect 16724 8812 16820 8828
rect 15731 8760 16453 8761
rect 15731 8040 15732 8760
rect 16452 8040 16453 8760
rect 15731 8039 16453 8040
rect 15312 7972 15408 7988
rect 16724 7988 16740 8812
rect 16804 7988 16820 8812
rect 18136 8812 18232 8828
rect 17143 8760 17865 8761
rect 17143 8040 17144 8760
rect 17864 8040 17865 8760
rect 17143 8039 17865 8040
rect 16724 7972 16820 7988
rect 18136 7988 18152 8812
rect 18216 7988 18232 8812
rect 19548 8812 19644 8828
rect 18555 8760 19277 8761
rect 18555 8040 18556 8760
rect 19276 8040 19277 8760
rect 18555 8039 19277 8040
rect 18136 7972 18232 7988
rect 19548 7988 19564 8812
rect 19628 7988 19644 8812
rect 20960 8812 21056 8828
rect 19967 8760 20689 8761
rect 19967 8040 19968 8760
rect 20688 8040 20689 8760
rect 19967 8039 20689 8040
rect 19548 7972 19644 7988
rect 20960 7988 20976 8812
rect 21040 7988 21056 8812
rect 22372 8812 22468 8828
rect 21379 8760 22101 8761
rect 21379 8040 21380 8760
rect 22100 8040 22101 8760
rect 21379 8039 22101 8040
rect 20960 7972 21056 7988
rect 22372 7988 22388 8812
rect 22452 7988 22468 8812
rect 23784 8812 23880 8828
rect 22791 8760 23513 8761
rect 22791 8040 22792 8760
rect 23512 8040 23513 8760
rect 22791 8039 23513 8040
rect 22372 7972 22468 7988
rect 23784 7988 23800 8812
rect 23864 7988 23880 8812
rect 23784 7972 23880 7988
rect -22812 7692 -22716 7708
rect -23805 7640 -23083 7641
rect -23805 6920 -23804 7640
rect -23084 6920 -23083 7640
rect -23805 6919 -23083 6920
rect -22812 6868 -22796 7692
rect -22732 6868 -22716 7692
rect -21400 7692 -21304 7708
rect -22393 7640 -21671 7641
rect -22393 6920 -22392 7640
rect -21672 6920 -21671 7640
rect -22393 6919 -21671 6920
rect -22812 6852 -22716 6868
rect -21400 6868 -21384 7692
rect -21320 6868 -21304 7692
rect -19988 7692 -19892 7708
rect -20981 7640 -20259 7641
rect -20981 6920 -20980 7640
rect -20260 6920 -20259 7640
rect -20981 6919 -20259 6920
rect -21400 6852 -21304 6868
rect -19988 6868 -19972 7692
rect -19908 6868 -19892 7692
rect -18576 7692 -18480 7708
rect -19569 7640 -18847 7641
rect -19569 6920 -19568 7640
rect -18848 6920 -18847 7640
rect -19569 6919 -18847 6920
rect -19988 6852 -19892 6868
rect -18576 6868 -18560 7692
rect -18496 6868 -18480 7692
rect -17164 7692 -17068 7708
rect -18157 7640 -17435 7641
rect -18157 6920 -18156 7640
rect -17436 6920 -17435 7640
rect -18157 6919 -17435 6920
rect -18576 6852 -18480 6868
rect -17164 6868 -17148 7692
rect -17084 6868 -17068 7692
rect -15752 7692 -15656 7708
rect -16745 7640 -16023 7641
rect -16745 6920 -16744 7640
rect -16024 6920 -16023 7640
rect -16745 6919 -16023 6920
rect -17164 6852 -17068 6868
rect -15752 6868 -15736 7692
rect -15672 6868 -15656 7692
rect -14340 7692 -14244 7708
rect -15333 7640 -14611 7641
rect -15333 6920 -15332 7640
rect -14612 6920 -14611 7640
rect -15333 6919 -14611 6920
rect -15752 6852 -15656 6868
rect -14340 6868 -14324 7692
rect -14260 6868 -14244 7692
rect -12928 7692 -12832 7708
rect -13921 7640 -13199 7641
rect -13921 6920 -13920 7640
rect -13200 6920 -13199 7640
rect -13921 6919 -13199 6920
rect -14340 6852 -14244 6868
rect -12928 6868 -12912 7692
rect -12848 6868 -12832 7692
rect -11516 7692 -11420 7708
rect -12509 7640 -11787 7641
rect -12509 6920 -12508 7640
rect -11788 6920 -11787 7640
rect -12509 6919 -11787 6920
rect -12928 6852 -12832 6868
rect -11516 6868 -11500 7692
rect -11436 6868 -11420 7692
rect -10104 7692 -10008 7708
rect -11097 7640 -10375 7641
rect -11097 6920 -11096 7640
rect -10376 6920 -10375 7640
rect -11097 6919 -10375 6920
rect -11516 6852 -11420 6868
rect -10104 6868 -10088 7692
rect -10024 6868 -10008 7692
rect -8692 7692 -8596 7708
rect -9685 7640 -8963 7641
rect -9685 6920 -9684 7640
rect -8964 6920 -8963 7640
rect -9685 6919 -8963 6920
rect -10104 6852 -10008 6868
rect -8692 6868 -8676 7692
rect -8612 6868 -8596 7692
rect -7280 7692 -7184 7708
rect -8273 7640 -7551 7641
rect -8273 6920 -8272 7640
rect -7552 6920 -7551 7640
rect -8273 6919 -7551 6920
rect -8692 6852 -8596 6868
rect -7280 6868 -7264 7692
rect -7200 6868 -7184 7692
rect -5868 7692 -5772 7708
rect -6861 7640 -6139 7641
rect -6861 6920 -6860 7640
rect -6140 6920 -6139 7640
rect -6861 6919 -6139 6920
rect -7280 6852 -7184 6868
rect -5868 6868 -5852 7692
rect -5788 6868 -5772 7692
rect -4456 7692 -4360 7708
rect -5449 7640 -4727 7641
rect -5449 6920 -5448 7640
rect -4728 6920 -4727 7640
rect -5449 6919 -4727 6920
rect -5868 6852 -5772 6868
rect -4456 6868 -4440 7692
rect -4376 6868 -4360 7692
rect -3044 7692 -2948 7708
rect -4037 7640 -3315 7641
rect -4037 6920 -4036 7640
rect -3316 6920 -3315 7640
rect -4037 6919 -3315 6920
rect -4456 6852 -4360 6868
rect -3044 6868 -3028 7692
rect -2964 6868 -2948 7692
rect -1632 7692 -1536 7708
rect -2625 7640 -1903 7641
rect -2625 6920 -2624 7640
rect -1904 6920 -1903 7640
rect -2625 6919 -1903 6920
rect -3044 6852 -2948 6868
rect -1632 6868 -1616 7692
rect -1552 6868 -1536 7692
rect -220 7692 -124 7708
rect -1213 7640 -491 7641
rect -1213 6920 -1212 7640
rect -492 6920 -491 7640
rect -1213 6919 -491 6920
rect -1632 6852 -1536 6868
rect -220 6868 -204 7692
rect -140 6868 -124 7692
rect 1192 7692 1288 7708
rect 199 7640 921 7641
rect 199 6920 200 7640
rect 920 6920 921 7640
rect 199 6919 921 6920
rect -220 6852 -124 6868
rect 1192 6868 1208 7692
rect 1272 6868 1288 7692
rect 2604 7692 2700 7708
rect 1611 7640 2333 7641
rect 1611 6920 1612 7640
rect 2332 6920 2333 7640
rect 1611 6919 2333 6920
rect 1192 6852 1288 6868
rect 2604 6868 2620 7692
rect 2684 6868 2700 7692
rect 4016 7692 4112 7708
rect 3023 7640 3745 7641
rect 3023 6920 3024 7640
rect 3744 6920 3745 7640
rect 3023 6919 3745 6920
rect 2604 6852 2700 6868
rect 4016 6868 4032 7692
rect 4096 6868 4112 7692
rect 5428 7692 5524 7708
rect 4435 7640 5157 7641
rect 4435 6920 4436 7640
rect 5156 6920 5157 7640
rect 4435 6919 5157 6920
rect 4016 6852 4112 6868
rect 5428 6868 5444 7692
rect 5508 6868 5524 7692
rect 6840 7692 6936 7708
rect 5847 7640 6569 7641
rect 5847 6920 5848 7640
rect 6568 6920 6569 7640
rect 5847 6919 6569 6920
rect 5428 6852 5524 6868
rect 6840 6868 6856 7692
rect 6920 6868 6936 7692
rect 8252 7692 8348 7708
rect 7259 7640 7981 7641
rect 7259 6920 7260 7640
rect 7980 6920 7981 7640
rect 7259 6919 7981 6920
rect 6840 6852 6936 6868
rect 8252 6868 8268 7692
rect 8332 6868 8348 7692
rect 9664 7692 9760 7708
rect 8671 7640 9393 7641
rect 8671 6920 8672 7640
rect 9392 6920 9393 7640
rect 8671 6919 9393 6920
rect 8252 6852 8348 6868
rect 9664 6868 9680 7692
rect 9744 6868 9760 7692
rect 11076 7692 11172 7708
rect 10083 7640 10805 7641
rect 10083 6920 10084 7640
rect 10804 6920 10805 7640
rect 10083 6919 10805 6920
rect 9664 6852 9760 6868
rect 11076 6868 11092 7692
rect 11156 6868 11172 7692
rect 12488 7692 12584 7708
rect 11495 7640 12217 7641
rect 11495 6920 11496 7640
rect 12216 6920 12217 7640
rect 11495 6919 12217 6920
rect 11076 6852 11172 6868
rect 12488 6868 12504 7692
rect 12568 6868 12584 7692
rect 13900 7692 13996 7708
rect 12907 7640 13629 7641
rect 12907 6920 12908 7640
rect 13628 6920 13629 7640
rect 12907 6919 13629 6920
rect 12488 6852 12584 6868
rect 13900 6868 13916 7692
rect 13980 6868 13996 7692
rect 15312 7692 15408 7708
rect 14319 7640 15041 7641
rect 14319 6920 14320 7640
rect 15040 6920 15041 7640
rect 14319 6919 15041 6920
rect 13900 6852 13996 6868
rect 15312 6868 15328 7692
rect 15392 6868 15408 7692
rect 16724 7692 16820 7708
rect 15731 7640 16453 7641
rect 15731 6920 15732 7640
rect 16452 6920 16453 7640
rect 15731 6919 16453 6920
rect 15312 6852 15408 6868
rect 16724 6868 16740 7692
rect 16804 6868 16820 7692
rect 18136 7692 18232 7708
rect 17143 7640 17865 7641
rect 17143 6920 17144 7640
rect 17864 6920 17865 7640
rect 17143 6919 17865 6920
rect 16724 6852 16820 6868
rect 18136 6868 18152 7692
rect 18216 6868 18232 7692
rect 19548 7692 19644 7708
rect 18555 7640 19277 7641
rect 18555 6920 18556 7640
rect 19276 6920 19277 7640
rect 18555 6919 19277 6920
rect 18136 6852 18232 6868
rect 19548 6868 19564 7692
rect 19628 6868 19644 7692
rect 20960 7692 21056 7708
rect 19967 7640 20689 7641
rect 19967 6920 19968 7640
rect 20688 6920 20689 7640
rect 19967 6919 20689 6920
rect 19548 6852 19644 6868
rect 20960 6868 20976 7692
rect 21040 6868 21056 7692
rect 22372 7692 22468 7708
rect 21379 7640 22101 7641
rect 21379 6920 21380 7640
rect 22100 6920 22101 7640
rect 21379 6919 22101 6920
rect 20960 6852 21056 6868
rect 22372 6868 22388 7692
rect 22452 6868 22468 7692
rect 23784 7692 23880 7708
rect 22791 7640 23513 7641
rect 22791 6920 22792 7640
rect 23512 6920 23513 7640
rect 22791 6919 23513 6920
rect 22372 6852 22468 6868
rect 23784 6868 23800 7692
rect 23864 6868 23880 7692
rect 23784 6852 23880 6868
rect -22812 6572 -22716 6588
rect -23805 6520 -23083 6521
rect -23805 5800 -23804 6520
rect -23084 5800 -23083 6520
rect -23805 5799 -23083 5800
rect -22812 5748 -22796 6572
rect -22732 5748 -22716 6572
rect -21400 6572 -21304 6588
rect -22393 6520 -21671 6521
rect -22393 5800 -22392 6520
rect -21672 5800 -21671 6520
rect -22393 5799 -21671 5800
rect -22812 5732 -22716 5748
rect -21400 5748 -21384 6572
rect -21320 5748 -21304 6572
rect -19988 6572 -19892 6588
rect -20981 6520 -20259 6521
rect -20981 5800 -20980 6520
rect -20260 5800 -20259 6520
rect -20981 5799 -20259 5800
rect -21400 5732 -21304 5748
rect -19988 5748 -19972 6572
rect -19908 5748 -19892 6572
rect -18576 6572 -18480 6588
rect -19569 6520 -18847 6521
rect -19569 5800 -19568 6520
rect -18848 5800 -18847 6520
rect -19569 5799 -18847 5800
rect -19988 5732 -19892 5748
rect -18576 5748 -18560 6572
rect -18496 5748 -18480 6572
rect -17164 6572 -17068 6588
rect -18157 6520 -17435 6521
rect -18157 5800 -18156 6520
rect -17436 5800 -17435 6520
rect -18157 5799 -17435 5800
rect -18576 5732 -18480 5748
rect -17164 5748 -17148 6572
rect -17084 5748 -17068 6572
rect -15752 6572 -15656 6588
rect -16745 6520 -16023 6521
rect -16745 5800 -16744 6520
rect -16024 5800 -16023 6520
rect -16745 5799 -16023 5800
rect -17164 5732 -17068 5748
rect -15752 5748 -15736 6572
rect -15672 5748 -15656 6572
rect -14340 6572 -14244 6588
rect -15333 6520 -14611 6521
rect -15333 5800 -15332 6520
rect -14612 5800 -14611 6520
rect -15333 5799 -14611 5800
rect -15752 5732 -15656 5748
rect -14340 5748 -14324 6572
rect -14260 5748 -14244 6572
rect -12928 6572 -12832 6588
rect -13921 6520 -13199 6521
rect -13921 5800 -13920 6520
rect -13200 5800 -13199 6520
rect -13921 5799 -13199 5800
rect -14340 5732 -14244 5748
rect -12928 5748 -12912 6572
rect -12848 5748 -12832 6572
rect -11516 6572 -11420 6588
rect -12509 6520 -11787 6521
rect -12509 5800 -12508 6520
rect -11788 5800 -11787 6520
rect -12509 5799 -11787 5800
rect -12928 5732 -12832 5748
rect -11516 5748 -11500 6572
rect -11436 5748 -11420 6572
rect -10104 6572 -10008 6588
rect -11097 6520 -10375 6521
rect -11097 5800 -11096 6520
rect -10376 5800 -10375 6520
rect -11097 5799 -10375 5800
rect -11516 5732 -11420 5748
rect -10104 5748 -10088 6572
rect -10024 5748 -10008 6572
rect -8692 6572 -8596 6588
rect -9685 6520 -8963 6521
rect -9685 5800 -9684 6520
rect -8964 5800 -8963 6520
rect -9685 5799 -8963 5800
rect -10104 5732 -10008 5748
rect -8692 5748 -8676 6572
rect -8612 5748 -8596 6572
rect -7280 6572 -7184 6588
rect -8273 6520 -7551 6521
rect -8273 5800 -8272 6520
rect -7552 5800 -7551 6520
rect -8273 5799 -7551 5800
rect -8692 5732 -8596 5748
rect -7280 5748 -7264 6572
rect -7200 5748 -7184 6572
rect -5868 6572 -5772 6588
rect -6861 6520 -6139 6521
rect -6861 5800 -6860 6520
rect -6140 5800 -6139 6520
rect -6861 5799 -6139 5800
rect -7280 5732 -7184 5748
rect -5868 5748 -5852 6572
rect -5788 5748 -5772 6572
rect -4456 6572 -4360 6588
rect -5449 6520 -4727 6521
rect -5449 5800 -5448 6520
rect -4728 5800 -4727 6520
rect -5449 5799 -4727 5800
rect -5868 5732 -5772 5748
rect -4456 5748 -4440 6572
rect -4376 5748 -4360 6572
rect -3044 6572 -2948 6588
rect -4037 6520 -3315 6521
rect -4037 5800 -4036 6520
rect -3316 5800 -3315 6520
rect -4037 5799 -3315 5800
rect -4456 5732 -4360 5748
rect -3044 5748 -3028 6572
rect -2964 5748 -2948 6572
rect -1632 6572 -1536 6588
rect -2625 6520 -1903 6521
rect -2625 5800 -2624 6520
rect -1904 5800 -1903 6520
rect -2625 5799 -1903 5800
rect -3044 5732 -2948 5748
rect -1632 5748 -1616 6572
rect -1552 5748 -1536 6572
rect -220 6572 -124 6588
rect -1213 6520 -491 6521
rect -1213 5800 -1212 6520
rect -492 5800 -491 6520
rect -1213 5799 -491 5800
rect -1632 5732 -1536 5748
rect -220 5748 -204 6572
rect -140 5748 -124 6572
rect 1192 6572 1288 6588
rect 199 6520 921 6521
rect 199 5800 200 6520
rect 920 5800 921 6520
rect 199 5799 921 5800
rect -220 5732 -124 5748
rect 1192 5748 1208 6572
rect 1272 5748 1288 6572
rect 2604 6572 2700 6588
rect 1611 6520 2333 6521
rect 1611 5800 1612 6520
rect 2332 5800 2333 6520
rect 1611 5799 2333 5800
rect 1192 5732 1288 5748
rect 2604 5748 2620 6572
rect 2684 5748 2700 6572
rect 4016 6572 4112 6588
rect 3023 6520 3745 6521
rect 3023 5800 3024 6520
rect 3744 5800 3745 6520
rect 3023 5799 3745 5800
rect 2604 5732 2700 5748
rect 4016 5748 4032 6572
rect 4096 5748 4112 6572
rect 5428 6572 5524 6588
rect 4435 6520 5157 6521
rect 4435 5800 4436 6520
rect 5156 5800 5157 6520
rect 4435 5799 5157 5800
rect 4016 5732 4112 5748
rect 5428 5748 5444 6572
rect 5508 5748 5524 6572
rect 6840 6572 6936 6588
rect 5847 6520 6569 6521
rect 5847 5800 5848 6520
rect 6568 5800 6569 6520
rect 5847 5799 6569 5800
rect 5428 5732 5524 5748
rect 6840 5748 6856 6572
rect 6920 5748 6936 6572
rect 8252 6572 8348 6588
rect 7259 6520 7981 6521
rect 7259 5800 7260 6520
rect 7980 5800 7981 6520
rect 7259 5799 7981 5800
rect 6840 5732 6936 5748
rect 8252 5748 8268 6572
rect 8332 5748 8348 6572
rect 9664 6572 9760 6588
rect 8671 6520 9393 6521
rect 8671 5800 8672 6520
rect 9392 5800 9393 6520
rect 8671 5799 9393 5800
rect 8252 5732 8348 5748
rect 9664 5748 9680 6572
rect 9744 5748 9760 6572
rect 11076 6572 11172 6588
rect 10083 6520 10805 6521
rect 10083 5800 10084 6520
rect 10804 5800 10805 6520
rect 10083 5799 10805 5800
rect 9664 5732 9760 5748
rect 11076 5748 11092 6572
rect 11156 5748 11172 6572
rect 12488 6572 12584 6588
rect 11495 6520 12217 6521
rect 11495 5800 11496 6520
rect 12216 5800 12217 6520
rect 11495 5799 12217 5800
rect 11076 5732 11172 5748
rect 12488 5748 12504 6572
rect 12568 5748 12584 6572
rect 13900 6572 13996 6588
rect 12907 6520 13629 6521
rect 12907 5800 12908 6520
rect 13628 5800 13629 6520
rect 12907 5799 13629 5800
rect 12488 5732 12584 5748
rect 13900 5748 13916 6572
rect 13980 5748 13996 6572
rect 15312 6572 15408 6588
rect 14319 6520 15041 6521
rect 14319 5800 14320 6520
rect 15040 5800 15041 6520
rect 14319 5799 15041 5800
rect 13900 5732 13996 5748
rect 15312 5748 15328 6572
rect 15392 5748 15408 6572
rect 16724 6572 16820 6588
rect 15731 6520 16453 6521
rect 15731 5800 15732 6520
rect 16452 5800 16453 6520
rect 15731 5799 16453 5800
rect 15312 5732 15408 5748
rect 16724 5748 16740 6572
rect 16804 5748 16820 6572
rect 18136 6572 18232 6588
rect 17143 6520 17865 6521
rect 17143 5800 17144 6520
rect 17864 5800 17865 6520
rect 17143 5799 17865 5800
rect 16724 5732 16820 5748
rect 18136 5748 18152 6572
rect 18216 5748 18232 6572
rect 19548 6572 19644 6588
rect 18555 6520 19277 6521
rect 18555 5800 18556 6520
rect 19276 5800 19277 6520
rect 18555 5799 19277 5800
rect 18136 5732 18232 5748
rect 19548 5748 19564 6572
rect 19628 5748 19644 6572
rect 20960 6572 21056 6588
rect 19967 6520 20689 6521
rect 19967 5800 19968 6520
rect 20688 5800 20689 6520
rect 19967 5799 20689 5800
rect 19548 5732 19644 5748
rect 20960 5748 20976 6572
rect 21040 5748 21056 6572
rect 22372 6572 22468 6588
rect 21379 6520 22101 6521
rect 21379 5800 21380 6520
rect 22100 5800 22101 6520
rect 21379 5799 22101 5800
rect 20960 5732 21056 5748
rect 22372 5748 22388 6572
rect 22452 5748 22468 6572
rect 23784 6572 23880 6588
rect 22791 6520 23513 6521
rect 22791 5800 22792 6520
rect 23512 5800 23513 6520
rect 22791 5799 23513 5800
rect 22372 5732 22468 5748
rect 23784 5748 23800 6572
rect 23864 5748 23880 6572
rect 23784 5732 23880 5748
rect -22812 5452 -22716 5468
rect -23805 5400 -23083 5401
rect -23805 4680 -23804 5400
rect -23084 4680 -23083 5400
rect -23805 4679 -23083 4680
rect -22812 4628 -22796 5452
rect -22732 4628 -22716 5452
rect -21400 5452 -21304 5468
rect -22393 5400 -21671 5401
rect -22393 4680 -22392 5400
rect -21672 4680 -21671 5400
rect -22393 4679 -21671 4680
rect -22812 4612 -22716 4628
rect -21400 4628 -21384 5452
rect -21320 4628 -21304 5452
rect -19988 5452 -19892 5468
rect -20981 5400 -20259 5401
rect -20981 4680 -20980 5400
rect -20260 4680 -20259 5400
rect -20981 4679 -20259 4680
rect -21400 4612 -21304 4628
rect -19988 4628 -19972 5452
rect -19908 4628 -19892 5452
rect -18576 5452 -18480 5468
rect -19569 5400 -18847 5401
rect -19569 4680 -19568 5400
rect -18848 4680 -18847 5400
rect -19569 4679 -18847 4680
rect -19988 4612 -19892 4628
rect -18576 4628 -18560 5452
rect -18496 4628 -18480 5452
rect -17164 5452 -17068 5468
rect -18157 5400 -17435 5401
rect -18157 4680 -18156 5400
rect -17436 4680 -17435 5400
rect -18157 4679 -17435 4680
rect -18576 4612 -18480 4628
rect -17164 4628 -17148 5452
rect -17084 4628 -17068 5452
rect -15752 5452 -15656 5468
rect -16745 5400 -16023 5401
rect -16745 4680 -16744 5400
rect -16024 4680 -16023 5400
rect -16745 4679 -16023 4680
rect -17164 4612 -17068 4628
rect -15752 4628 -15736 5452
rect -15672 4628 -15656 5452
rect -14340 5452 -14244 5468
rect -15333 5400 -14611 5401
rect -15333 4680 -15332 5400
rect -14612 4680 -14611 5400
rect -15333 4679 -14611 4680
rect -15752 4612 -15656 4628
rect -14340 4628 -14324 5452
rect -14260 4628 -14244 5452
rect -12928 5452 -12832 5468
rect -13921 5400 -13199 5401
rect -13921 4680 -13920 5400
rect -13200 4680 -13199 5400
rect -13921 4679 -13199 4680
rect -14340 4612 -14244 4628
rect -12928 4628 -12912 5452
rect -12848 4628 -12832 5452
rect -11516 5452 -11420 5468
rect -12509 5400 -11787 5401
rect -12509 4680 -12508 5400
rect -11788 4680 -11787 5400
rect -12509 4679 -11787 4680
rect -12928 4612 -12832 4628
rect -11516 4628 -11500 5452
rect -11436 4628 -11420 5452
rect -10104 5452 -10008 5468
rect -11097 5400 -10375 5401
rect -11097 4680 -11096 5400
rect -10376 4680 -10375 5400
rect -11097 4679 -10375 4680
rect -11516 4612 -11420 4628
rect -10104 4628 -10088 5452
rect -10024 4628 -10008 5452
rect -8692 5452 -8596 5468
rect -9685 5400 -8963 5401
rect -9685 4680 -9684 5400
rect -8964 4680 -8963 5400
rect -9685 4679 -8963 4680
rect -10104 4612 -10008 4628
rect -8692 4628 -8676 5452
rect -8612 4628 -8596 5452
rect -7280 5452 -7184 5468
rect -8273 5400 -7551 5401
rect -8273 4680 -8272 5400
rect -7552 4680 -7551 5400
rect -8273 4679 -7551 4680
rect -8692 4612 -8596 4628
rect -7280 4628 -7264 5452
rect -7200 4628 -7184 5452
rect -5868 5452 -5772 5468
rect -6861 5400 -6139 5401
rect -6861 4680 -6860 5400
rect -6140 4680 -6139 5400
rect -6861 4679 -6139 4680
rect -7280 4612 -7184 4628
rect -5868 4628 -5852 5452
rect -5788 4628 -5772 5452
rect -4456 5452 -4360 5468
rect -5449 5400 -4727 5401
rect -5449 4680 -5448 5400
rect -4728 4680 -4727 5400
rect -5449 4679 -4727 4680
rect -5868 4612 -5772 4628
rect -4456 4628 -4440 5452
rect -4376 4628 -4360 5452
rect -3044 5452 -2948 5468
rect -4037 5400 -3315 5401
rect -4037 4680 -4036 5400
rect -3316 4680 -3315 5400
rect -4037 4679 -3315 4680
rect -4456 4612 -4360 4628
rect -3044 4628 -3028 5452
rect -2964 4628 -2948 5452
rect -1632 5452 -1536 5468
rect -2625 5400 -1903 5401
rect -2625 4680 -2624 5400
rect -1904 4680 -1903 5400
rect -2625 4679 -1903 4680
rect -3044 4612 -2948 4628
rect -1632 4628 -1616 5452
rect -1552 4628 -1536 5452
rect -220 5452 -124 5468
rect -1213 5400 -491 5401
rect -1213 4680 -1212 5400
rect -492 4680 -491 5400
rect -1213 4679 -491 4680
rect -1632 4612 -1536 4628
rect -220 4628 -204 5452
rect -140 4628 -124 5452
rect 1192 5452 1288 5468
rect 199 5400 921 5401
rect 199 4680 200 5400
rect 920 4680 921 5400
rect 199 4679 921 4680
rect -220 4612 -124 4628
rect 1192 4628 1208 5452
rect 1272 4628 1288 5452
rect 2604 5452 2700 5468
rect 1611 5400 2333 5401
rect 1611 4680 1612 5400
rect 2332 4680 2333 5400
rect 1611 4679 2333 4680
rect 1192 4612 1288 4628
rect 2604 4628 2620 5452
rect 2684 4628 2700 5452
rect 4016 5452 4112 5468
rect 3023 5400 3745 5401
rect 3023 4680 3024 5400
rect 3744 4680 3745 5400
rect 3023 4679 3745 4680
rect 2604 4612 2700 4628
rect 4016 4628 4032 5452
rect 4096 4628 4112 5452
rect 5428 5452 5524 5468
rect 4435 5400 5157 5401
rect 4435 4680 4436 5400
rect 5156 4680 5157 5400
rect 4435 4679 5157 4680
rect 4016 4612 4112 4628
rect 5428 4628 5444 5452
rect 5508 4628 5524 5452
rect 6840 5452 6936 5468
rect 5847 5400 6569 5401
rect 5847 4680 5848 5400
rect 6568 4680 6569 5400
rect 5847 4679 6569 4680
rect 5428 4612 5524 4628
rect 6840 4628 6856 5452
rect 6920 4628 6936 5452
rect 8252 5452 8348 5468
rect 7259 5400 7981 5401
rect 7259 4680 7260 5400
rect 7980 4680 7981 5400
rect 7259 4679 7981 4680
rect 6840 4612 6936 4628
rect 8252 4628 8268 5452
rect 8332 4628 8348 5452
rect 9664 5452 9760 5468
rect 8671 5400 9393 5401
rect 8671 4680 8672 5400
rect 9392 4680 9393 5400
rect 8671 4679 9393 4680
rect 8252 4612 8348 4628
rect 9664 4628 9680 5452
rect 9744 4628 9760 5452
rect 11076 5452 11172 5468
rect 10083 5400 10805 5401
rect 10083 4680 10084 5400
rect 10804 4680 10805 5400
rect 10083 4679 10805 4680
rect 9664 4612 9760 4628
rect 11076 4628 11092 5452
rect 11156 4628 11172 5452
rect 12488 5452 12584 5468
rect 11495 5400 12217 5401
rect 11495 4680 11496 5400
rect 12216 4680 12217 5400
rect 11495 4679 12217 4680
rect 11076 4612 11172 4628
rect 12488 4628 12504 5452
rect 12568 4628 12584 5452
rect 13900 5452 13996 5468
rect 12907 5400 13629 5401
rect 12907 4680 12908 5400
rect 13628 4680 13629 5400
rect 12907 4679 13629 4680
rect 12488 4612 12584 4628
rect 13900 4628 13916 5452
rect 13980 4628 13996 5452
rect 15312 5452 15408 5468
rect 14319 5400 15041 5401
rect 14319 4680 14320 5400
rect 15040 4680 15041 5400
rect 14319 4679 15041 4680
rect 13900 4612 13996 4628
rect 15312 4628 15328 5452
rect 15392 4628 15408 5452
rect 16724 5452 16820 5468
rect 15731 5400 16453 5401
rect 15731 4680 15732 5400
rect 16452 4680 16453 5400
rect 15731 4679 16453 4680
rect 15312 4612 15408 4628
rect 16724 4628 16740 5452
rect 16804 4628 16820 5452
rect 18136 5452 18232 5468
rect 17143 5400 17865 5401
rect 17143 4680 17144 5400
rect 17864 4680 17865 5400
rect 17143 4679 17865 4680
rect 16724 4612 16820 4628
rect 18136 4628 18152 5452
rect 18216 4628 18232 5452
rect 19548 5452 19644 5468
rect 18555 5400 19277 5401
rect 18555 4680 18556 5400
rect 19276 4680 19277 5400
rect 18555 4679 19277 4680
rect 18136 4612 18232 4628
rect 19548 4628 19564 5452
rect 19628 4628 19644 5452
rect 20960 5452 21056 5468
rect 19967 5400 20689 5401
rect 19967 4680 19968 5400
rect 20688 4680 20689 5400
rect 19967 4679 20689 4680
rect 19548 4612 19644 4628
rect 20960 4628 20976 5452
rect 21040 4628 21056 5452
rect 22372 5452 22468 5468
rect 21379 5400 22101 5401
rect 21379 4680 21380 5400
rect 22100 4680 22101 5400
rect 21379 4679 22101 4680
rect 20960 4612 21056 4628
rect 22372 4628 22388 5452
rect 22452 4628 22468 5452
rect 23784 5452 23880 5468
rect 22791 5400 23513 5401
rect 22791 4680 22792 5400
rect 23512 4680 23513 5400
rect 22791 4679 23513 4680
rect 22372 4612 22468 4628
rect 23784 4628 23800 5452
rect 23864 4628 23880 5452
rect 23784 4612 23880 4628
rect -22812 4332 -22716 4348
rect -23805 4280 -23083 4281
rect -23805 3560 -23804 4280
rect -23084 3560 -23083 4280
rect -23805 3559 -23083 3560
rect -22812 3508 -22796 4332
rect -22732 3508 -22716 4332
rect -21400 4332 -21304 4348
rect -22393 4280 -21671 4281
rect -22393 3560 -22392 4280
rect -21672 3560 -21671 4280
rect -22393 3559 -21671 3560
rect -22812 3492 -22716 3508
rect -21400 3508 -21384 4332
rect -21320 3508 -21304 4332
rect -19988 4332 -19892 4348
rect -20981 4280 -20259 4281
rect -20981 3560 -20980 4280
rect -20260 3560 -20259 4280
rect -20981 3559 -20259 3560
rect -21400 3492 -21304 3508
rect -19988 3508 -19972 4332
rect -19908 3508 -19892 4332
rect -18576 4332 -18480 4348
rect -19569 4280 -18847 4281
rect -19569 3560 -19568 4280
rect -18848 3560 -18847 4280
rect -19569 3559 -18847 3560
rect -19988 3492 -19892 3508
rect -18576 3508 -18560 4332
rect -18496 3508 -18480 4332
rect -17164 4332 -17068 4348
rect -18157 4280 -17435 4281
rect -18157 3560 -18156 4280
rect -17436 3560 -17435 4280
rect -18157 3559 -17435 3560
rect -18576 3492 -18480 3508
rect -17164 3508 -17148 4332
rect -17084 3508 -17068 4332
rect -15752 4332 -15656 4348
rect -16745 4280 -16023 4281
rect -16745 3560 -16744 4280
rect -16024 3560 -16023 4280
rect -16745 3559 -16023 3560
rect -17164 3492 -17068 3508
rect -15752 3508 -15736 4332
rect -15672 3508 -15656 4332
rect -14340 4332 -14244 4348
rect -15333 4280 -14611 4281
rect -15333 3560 -15332 4280
rect -14612 3560 -14611 4280
rect -15333 3559 -14611 3560
rect -15752 3492 -15656 3508
rect -14340 3508 -14324 4332
rect -14260 3508 -14244 4332
rect -12928 4332 -12832 4348
rect -13921 4280 -13199 4281
rect -13921 3560 -13920 4280
rect -13200 3560 -13199 4280
rect -13921 3559 -13199 3560
rect -14340 3492 -14244 3508
rect -12928 3508 -12912 4332
rect -12848 3508 -12832 4332
rect -11516 4332 -11420 4348
rect -12509 4280 -11787 4281
rect -12509 3560 -12508 4280
rect -11788 3560 -11787 4280
rect -12509 3559 -11787 3560
rect -12928 3492 -12832 3508
rect -11516 3508 -11500 4332
rect -11436 3508 -11420 4332
rect -10104 4332 -10008 4348
rect -11097 4280 -10375 4281
rect -11097 3560 -11096 4280
rect -10376 3560 -10375 4280
rect -11097 3559 -10375 3560
rect -11516 3492 -11420 3508
rect -10104 3508 -10088 4332
rect -10024 3508 -10008 4332
rect -8692 4332 -8596 4348
rect -9685 4280 -8963 4281
rect -9685 3560 -9684 4280
rect -8964 3560 -8963 4280
rect -9685 3559 -8963 3560
rect -10104 3492 -10008 3508
rect -8692 3508 -8676 4332
rect -8612 3508 -8596 4332
rect -7280 4332 -7184 4348
rect -8273 4280 -7551 4281
rect -8273 3560 -8272 4280
rect -7552 3560 -7551 4280
rect -8273 3559 -7551 3560
rect -8692 3492 -8596 3508
rect -7280 3508 -7264 4332
rect -7200 3508 -7184 4332
rect -5868 4332 -5772 4348
rect -6861 4280 -6139 4281
rect -6861 3560 -6860 4280
rect -6140 3560 -6139 4280
rect -6861 3559 -6139 3560
rect -7280 3492 -7184 3508
rect -5868 3508 -5852 4332
rect -5788 3508 -5772 4332
rect -4456 4332 -4360 4348
rect -5449 4280 -4727 4281
rect -5449 3560 -5448 4280
rect -4728 3560 -4727 4280
rect -5449 3559 -4727 3560
rect -5868 3492 -5772 3508
rect -4456 3508 -4440 4332
rect -4376 3508 -4360 4332
rect -3044 4332 -2948 4348
rect -4037 4280 -3315 4281
rect -4037 3560 -4036 4280
rect -3316 3560 -3315 4280
rect -4037 3559 -3315 3560
rect -4456 3492 -4360 3508
rect -3044 3508 -3028 4332
rect -2964 3508 -2948 4332
rect -1632 4332 -1536 4348
rect -2625 4280 -1903 4281
rect -2625 3560 -2624 4280
rect -1904 3560 -1903 4280
rect -2625 3559 -1903 3560
rect -3044 3492 -2948 3508
rect -1632 3508 -1616 4332
rect -1552 3508 -1536 4332
rect -220 4332 -124 4348
rect -1213 4280 -491 4281
rect -1213 3560 -1212 4280
rect -492 3560 -491 4280
rect -1213 3559 -491 3560
rect -1632 3492 -1536 3508
rect -220 3508 -204 4332
rect -140 3508 -124 4332
rect 1192 4332 1288 4348
rect 199 4280 921 4281
rect 199 3560 200 4280
rect 920 3560 921 4280
rect 199 3559 921 3560
rect -220 3492 -124 3508
rect 1192 3508 1208 4332
rect 1272 3508 1288 4332
rect 2604 4332 2700 4348
rect 1611 4280 2333 4281
rect 1611 3560 1612 4280
rect 2332 3560 2333 4280
rect 1611 3559 2333 3560
rect 1192 3492 1288 3508
rect 2604 3508 2620 4332
rect 2684 3508 2700 4332
rect 4016 4332 4112 4348
rect 3023 4280 3745 4281
rect 3023 3560 3024 4280
rect 3744 3560 3745 4280
rect 3023 3559 3745 3560
rect 2604 3492 2700 3508
rect 4016 3508 4032 4332
rect 4096 3508 4112 4332
rect 5428 4332 5524 4348
rect 4435 4280 5157 4281
rect 4435 3560 4436 4280
rect 5156 3560 5157 4280
rect 4435 3559 5157 3560
rect 4016 3492 4112 3508
rect 5428 3508 5444 4332
rect 5508 3508 5524 4332
rect 6840 4332 6936 4348
rect 5847 4280 6569 4281
rect 5847 3560 5848 4280
rect 6568 3560 6569 4280
rect 5847 3559 6569 3560
rect 5428 3492 5524 3508
rect 6840 3508 6856 4332
rect 6920 3508 6936 4332
rect 8252 4332 8348 4348
rect 7259 4280 7981 4281
rect 7259 3560 7260 4280
rect 7980 3560 7981 4280
rect 7259 3559 7981 3560
rect 6840 3492 6936 3508
rect 8252 3508 8268 4332
rect 8332 3508 8348 4332
rect 9664 4332 9760 4348
rect 8671 4280 9393 4281
rect 8671 3560 8672 4280
rect 9392 3560 9393 4280
rect 8671 3559 9393 3560
rect 8252 3492 8348 3508
rect 9664 3508 9680 4332
rect 9744 3508 9760 4332
rect 11076 4332 11172 4348
rect 10083 4280 10805 4281
rect 10083 3560 10084 4280
rect 10804 3560 10805 4280
rect 10083 3559 10805 3560
rect 9664 3492 9760 3508
rect 11076 3508 11092 4332
rect 11156 3508 11172 4332
rect 12488 4332 12584 4348
rect 11495 4280 12217 4281
rect 11495 3560 11496 4280
rect 12216 3560 12217 4280
rect 11495 3559 12217 3560
rect 11076 3492 11172 3508
rect 12488 3508 12504 4332
rect 12568 3508 12584 4332
rect 13900 4332 13996 4348
rect 12907 4280 13629 4281
rect 12907 3560 12908 4280
rect 13628 3560 13629 4280
rect 12907 3559 13629 3560
rect 12488 3492 12584 3508
rect 13900 3508 13916 4332
rect 13980 3508 13996 4332
rect 15312 4332 15408 4348
rect 14319 4280 15041 4281
rect 14319 3560 14320 4280
rect 15040 3560 15041 4280
rect 14319 3559 15041 3560
rect 13900 3492 13996 3508
rect 15312 3508 15328 4332
rect 15392 3508 15408 4332
rect 16724 4332 16820 4348
rect 15731 4280 16453 4281
rect 15731 3560 15732 4280
rect 16452 3560 16453 4280
rect 15731 3559 16453 3560
rect 15312 3492 15408 3508
rect 16724 3508 16740 4332
rect 16804 3508 16820 4332
rect 18136 4332 18232 4348
rect 17143 4280 17865 4281
rect 17143 3560 17144 4280
rect 17864 3560 17865 4280
rect 17143 3559 17865 3560
rect 16724 3492 16820 3508
rect 18136 3508 18152 4332
rect 18216 3508 18232 4332
rect 19548 4332 19644 4348
rect 18555 4280 19277 4281
rect 18555 3560 18556 4280
rect 19276 3560 19277 4280
rect 18555 3559 19277 3560
rect 18136 3492 18232 3508
rect 19548 3508 19564 4332
rect 19628 3508 19644 4332
rect 20960 4332 21056 4348
rect 19967 4280 20689 4281
rect 19967 3560 19968 4280
rect 20688 3560 20689 4280
rect 19967 3559 20689 3560
rect 19548 3492 19644 3508
rect 20960 3508 20976 4332
rect 21040 3508 21056 4332
rect 22372 4332 22468 4348
rect 21379 4280 22101 4281
rect 21379 3560 21380 4280
rect 22100 3560 22101 4280
rect 21379 3559 22101 3560
rect 20960 3492 21056 3508
rect 22372 3508 22388 4332
rect 22452 3508 22468 4332
rect 23784 4332 23880 4348
rect 22791 4280 23513 4281
rect 22791 3560 22792 4280
rect 23512 3560 23513 4280
rect 22791 3559 23513 3560
rect 22372 3492 22468 3508
rect 23784 3508 23800 4332
rect 23864 3508 23880 4332
rect 23784 3492 23880 3508
rect -22812 3212 -22716 3228
rect -23805 3160 -23083 3161
rect -23805 2440 -23804 3160
rect -23084 2440 -23083 3160
rect -23805 2439 -23083 2440
rect -22812 2388 -22796 3212
rect -22732 2388 -22716 3212
rect -21400 3212 -21304 3228
rect -22393 3160 -21671 3161
rect -22393 2440 -22392 3160
rect -21672 2440 -21671 3160
rect -22393 2439 -21671 2440
rect -22812 2372 -22716 2388
rect -21400 2388 -21384 3212
rect -21320 2388 -21304 3212
rect -19988 3212 -19892 3228
rect -20981 3160 -20259 3161
rect -20981 2440 -20980 3160
rect -20260 2440 -20259 3160
rect -20981 2439 -20259 2440
rect -21400 2372 -21304 2388
rect -19988 2388 -19972 3212
rect -19908 2388 -19892 3212
rect -18576 3212 -18480 3228
rect -19569 3160 -18847 3161
rect -19569 2440 -19568 3160
rect -18848 2440 -18847 3160
rect -19569 2439 -18847 2440
rect -19988 2372 -19892 2388
rect -18576 2388 -18560 3212
rect -18496 2388 -18480 3212
rect -17164 3212 -17068 3228
rect -18157 3160 -17435 3161
rect -18157 2440 -18156 3160
rect -17436 2440 -17435 3160
rect -18157 2439 -17435 2440
rect -18576 2372 -18480 2388
rect -17164 2388 -17148 3212
rect -17084 2388 -17068 3212
rect -15752 3212 -15656 3228
rect -16745 3160 -16023 3161
rect -16745 2440 -16744 3160
rect -16024 2440 -16023 3160
rect -16745 2439 -16023 2440
rect -17164 2372 -17068 2388
rect -15752 2388 -15736 3212
rect -15672 2388 -15656 3212
rect -14340 3212 -14244 3228
rect -15333 3160 -14611 3161
rect -15333 2440 -15332 3160
rect -14612 2440 -14611 3160
rect -15333 2439 -14611 2440
rect -15752 2372 -15656 2388
rect -14340 2388 -14324 3212
rect -14260 2388 -14244 3212
rect -12928 3212 -12832 3228
rect -13921 3160 -13199 3161
rect -13921 2440 -13920 3160
rect -13200 2440 -13199 3160
rect -13921 2439 -13199 2440
rect -14340 2372 -14244 2388
rect -12928 2388 -12912 3212
rect -12848 2388 -12832 3212
rect -11516 3212 -11420 3228
rect -12509 3160 -11787 3161
rect -12509 2440 -12508 3160
rect -11788 2440 -11787 3160
rect -12509 2439 -11787 2440
rect -12928 2372 -12832 2388
rect -11516 2388 -11500 3212
rect -11436 2388 -11420 3212
rect -10104 3212 -10008 3228
rect -11097 3160 -10375 3161
rect -11097 2440 -11096 3160
rect -10376 2440 -10375 3160
rect -11097 2439 -10375 2440
rect -11516 2372 -11420 2388
rect -10104 2388 -10088 3212
rect -10024 2388 -10008 3212
rect -8692 3212 -8596 3228
rect -9685 3160 -8963 3161
rect -9685 2440 -9684 3160
rect -8964 2440 -8963 3160
rect -9685 2439 -8963 2440
rect -10104 2372 -10008 2388
rect -8692 2388 -8676 3212
rect -8612 2388 -8596 3212
rect -7280 3212 -7184 3228
rect -8273 3160 -7551 3161
rect -8273 2440 -8272 3160
rect -7552 2440 -7551 3160
rect -8273 2439 -7551 2440
rect -8692 2372 -8596 2388
rect -7280 2388 -7264 3212
rect -7200 2388 -7184 3212
rect -5868 3212 -5772 3228
rect -6861 3160 -6139 3161
rect -6861 2440 -6860 3160
rect -6140 2440 -6139 3160
rect -6861 2439 -6139 2440
rect -7280 2372 -7184 2388
rect -5868 2388 -5852 3212
rect -5788 2388 -5772 3212
rect -4456 3212 -4360 3228
rect -5449 3160 -4727 3161
rect -5449 2440 -5448 3160
rect -4728 2440 -4727 3160
rect -5449 2439 -4727 2440
rect -5868 2372 -5772 2388
rect -4456 2388 -4440 3212
rect -4376 2388 -4360 3212
rect -3044 3212 -2948 3228
rect -4037 3160 -3315 3161
rect -4037 2440 -4036 3160
rect -3316 2440 -3315 3160
rect -4037 2439 -3315 2440
rect -4456 2372 -4360 2388
rect -3044 2388 -3028 3212
rect -2964 2388 -2948 3212
rect -1632 3212 -1536 3228
rect -2625 3160 -1903 3161
rect -2625 2440 -2624 3160
rect -1904 2440 -1903 3160
rect -2625 2439 -1903 2440
rect -3044 2372 -2948 2388
rect -1632 2388 -1616 3212
rect -1552 2388 -1536 3212
rect -220 3212 -124 3228
rect -1213 3160 -491 3161
rect -1213 2440 -1212 3160
rect -492 2440 -491 3160
rect -1213 2439 -491 2440
rect -1632 2372 -1536 2388
rect -220 2388 -204 3212
rect -140 2388 -124 3212
rect 1192 3212 1288 3228
rect 199 3160 921 3161
rect 199 2440 200 3160
rect 920 2440 921 3160
rect 199 2439 921 2440
rect -220 2372 -124 2388
rect 1192 2388 1208 3212
rect 1272 2388 1288 3212
rect 2604 3212 2700 3228
rect 1611 3160 2333 3161
rect 1611 2440 1612 3160
rect 2332 2440 2333 3160
rect 1611 2439 2333 2440
rect 1192 2372 1288 2388
rect 2604 2388 2620 3212
rect 2684 2388 2700 3212
rect 4016 3212 4112 3228
rect 3023 3160 3745 3161
rect 3023 2440 3024 3160
rect 3744 2440 3745 3160
rect 3023 2439 3745 2440
rect 2604 2372 2700 2388
rect 4016 2388 4032 3212
rect 4096 2388 4112 3212
rect 5428 3212 5524 3228
rect 4435 3160 5157 3161
rect 4435 2440 4436 3160
rect 5156 2440 5157 3160
rect 4435 2439 5157 2440
rect 4016 2372 4112 2388
rect 5428 2388 5444 3212
rect 5508 2388 5524 3212
rect 6840 3212 6936 3228
rect 5847 3160 6569 3161
rect 5847 2440 5848 3160
rect 6568 2440 6569 3160
rect 5847 2439 6569 2440
rect 5428 2372 5524 2388
rect 6840 2388 6856 3212
rect 6920 2388 6936 3212
rect 8252 3212 8348 3228
rect 7259 3160 7981 3161
rect 7259 2440 7260 3160
rect 7980 2440 7981 3160
rect 7259 2439 7981 2440
rect 6840 2372 6936 2388
rect 8252 2388 8268 3212
rect 8332 2388 8348 3212
rect 9664 3212 9760 3228
rect 8671 3160 9393 3161
rect 8671 2440 8672 3160
rect 9392 2440 9393 3160
rect 8671 2439 9393 2440
rect 8252 2372 8348 2388
rect 9664 2388 9680 3212
rect 9744 2388 9760 3212
rect 11076 3212 11172 3228
rect 10083 3160 10805 3161
rect 10083 2440 10084 3160
rect 10804 2440 10805 3160
rect 10083 2439 10805 2440
rect 9664 2372 9760 2388
rect 11076 2388 11092 3212
rect 11156 2388 11172 3212
rect 12488 3212 12584 3228
rect 11495 3160 12217 3161
rect 11495 2440 11496 3160
rect 12216 2440 12217 3160
rect 11495 2439 12217 2440
rect 11076 2372 11172 2388
rect 12488 2388 12504 3212
rect 12568 2388 12584 3212
rect 13900 3212 13996 3228
rect 12907 3160 13629 3161
rect 12907 2440 12908 3160
rect 13628 2440 13629 3160
rect 12907 2439 13629 2440
rect 12488 2372 12584 2388
rect 13900 2388 13916 3212
rect 13980 2388 13996 3212
rect 15312 3212 15408 3228
rect 14319 3160 15041 3161
rect 14319 2440 14320 3160
rect 15040 2440 15041 3160
rect 14319 2439 15041 2440
rect 13900 2372 13996 2388
rect 15312 2388 15328 3212
rect 15392 2388 15408 3212
rect 16724 3212 16820 3228
rect 15731 3160 16453 3161
rect 15731 2440 15732 3160
rect 16452 2440 16453 3160
rect 15731 2439 16453 2440
rect 15312 2372 15408 2388
rect 16724 2388 16740 3212
rect 16804 2388 16820 3212
rect 18136 3212 18232 3228
rect 17143 3160 17865 3161
rect 17143 2440 17144 3160
rect 17864 2440 17865 3160
rect 17143 2439 17865 2440
rect 16724 2372 16820 2388
rect 18136 2388 18152 3212
rect 18216 2388 18232 3212
rect 19548 3212 19644 3228
rect 18555 3160 19277 3161
rect 18555 2440 18556 3160
rect 19276 2440 19277 3160
rect 18555 2439 19277 2440
rect 18136 2372 18232 2388
rect 19548 2388 19564 3212
rect 19628 2388 19644 3212
rect 20960 3212 21056 3228
rect 19967 3160 20689 3161
rect 19967 2440 19968 3160
rect 20688 2440 20689 3160
rect 19967 2439 20689 2440
rect 19548 2372 19644 2388
rect 20960 2388 20976 3212
rect 21040 2388 21056 3212
rect 22372 3212 22468 3228
rect 21379 3160 22101 3161
rect 21379 2440 21380 3160
rect 22100 2440 22101 3160
rect 21379 2439 22101 2440
rect 20960 2372 21056 2388
rect 22372 2388 22388 3212
rect 22452 2388 22468 3212
rect 23784 3212 23880 3228
rect 22791 3160 23513 3161
rect 22791 2440 22792 3160
rect 23512 2440 23513 3160
rect 22791 2439 23513 2440
rect 22372 2372 22468 2388
rect 23784 2388 23800 3212
rect 23864 2388 23880 3212
rect 23784 2372 23880 2388
rect -22812 2092 -22716 2108
rect -23805 2040 -23083 2041
rect -23805 1320 -23804 2040
rect -23084 1320 -23083 2040
rect -23805 1319 -23083 1320
rect -22812 1268 -22796 2092
rect -22732 1268 -22716 2092
rect -21400 2092 -21304 2108
rect -22393 2040 -21671 2041
rect -22393 1320 -22392 2040
rect -21672 1320 -21671 2040
rect -22393 1319 -21671 1320
rect -22812 1252 -22716 1268
rect -21400 1268 -21384 2092
rect -21320 1268 -21304 2092
rect -19988 2092 -19892 2108
rect -20981 2040 -20259 2041
rect -20981 1320 -20980 2040
rect -20260 1320 -20259 2040
rect -20981 1319 -20259 1320
rect -21400 1252 -21304 1268
rect -19988 1268 -19972 2092
rect -19908 1268 -19892 2092
rect -18576 2092 -18480 2108
rect -19569 2040 -18847 2041
rect -19569 1320 -19568 2040
rect -18848 1320 -18847 2040
rect -19569 1319 -18847 1320
rect -19988 1252 -19892 1268
rect -18576 1268 -18560 2092
rect -18496 1268 -18480 2092
rect -17164 2092 -17068 2108
rect -18157 2040 -17435 2041
rect -18157 1320 -18156 2040
rect -17436 1320 -17435 2040
rect -18157 1319 -17435 1320
rect -18576 1252 -18480 1268
rect -17164 1268 -17148 2092
rect -17084 1268 -17068 2092
rect -15752 2092 -15656 2108
rect -16745 2040 -16023 2041
rect -16745 1320 -16744 2040
rect -16024 1320 -16023 2040
rect -16745 1319 -16023 1320
rect -17164 1252 -17068 1268
rect -15752 1268 -15736 2092
rect -15672 1268 -15656 2092
rect -14340 2092 -14244 2108
rect -15333 2040 -14611 2041
rect -15333 1320 -15332 2040
rect -14612 1320 -14611 2040
rect -15333 1319 -14611 1320
rect -15752 1252 -15656 1268
rect -14340 1268 -14324 2092
rect -14260 1268 -14244 2092
rect -12928 2092 -12832 2108
rect -13921 2040 -13199 2041
rect -13921 1320 -13920 2040
rect -13200 1320 -13199 2040
rect -13921 1319 -13199 1320
rect -14340 1252 -14244 1268
rect -12928 1268 -12912 2092
rect -12848 1268 -12832 2092
rect -11516 2092 -11420 2108
rect -12509 2040 -11787 2041
rect -12509 1320 -12508 2040
rect -11788 1320 -11787 2040
rect -12509 1319 -11787 1320
rect -12928 1252 -12832 1268
rect -11516 1268 -11500 2092
rect -11436 1268 -11420 2092
rect -10104 2092 -10008 2108
rect -11097 2040 -10375 2041
rect -11097 1320 -11096 2040
rect -10376 1320 -10375 2040
rect -11097 1319 -10375 1320
rect -11516 1252 -11420 1268
rect -10104 1268 -10088 2092
rect -10024 1268 -10008 2092
rect -8692 2092 -8596 2108
rect -9685 2040 -8963 2041
rect -9685 1320 -9684 2040
rect -8964 1320 -8963 2040
rect -9685 1319 -8963 1320
rect -10104 1252 -10008 1268
rect -8692 1268 -8676 2092
rect -8612 1268 -8596 2092
rect -7280 2092 -7184 2108
rect -8273 2040 -7551 2041
rect -8273 1320 -8272 2040
rect -7552 1320 -7551 2040
rect -8273 1319 -7551 1320
rect -8692 1252 -8596 1268
rect -7280 1268 -7264 2092
rect -7200 1268 -7184 2092
rect -5868 2092 -5772 2108
rect -6861 2040 -6139 2041
rect -6861 1320 -6860 2040
rect -6140 1320 -6139 2040
rect -6861 1319 -6139 1320
rect -7280 1252 -7184 1268
rect -5868 1268 -5852 2092
rect -5788 1268 -5772 2092
rect -4456 2092 -4360 2108
rect -5449 2040 -4727 2041
rect -5449 1320 -5448 2040
rect -4728 1320 -4727 2040
rect -5449 1319 -4727 1320
rect -5868 1252 -5772 1268
rect -4456 1268 -4440 2092
rect -4376 1268 -4360 2092
rect -3044 2092 -2948 2108
rect -4037 2040 -3315 2041
rect -4037 1320 -4036 2040
rect -3316 1320 -3315 2040
rect -4037 1319 -3315 1320
rect -4456 1252 -4360 1268
rect -3044 1268 -3028 2092
rect -2964 1268 -2948 2092
rect -1632 2092 -1536 2108
rect -2625 2040 -1903 2041
rect -2625 1320 -2624 2040
rect -1904 1320 -1903 2040
rect -2625 1319 -1903 1320
rect -3044 1252 -2948 1268
rect -1632 1268 -1616 2092
rect -1552 1268 -1536 2092
rect -220 2092 -124 2108
rect -1213 2040 -491 2041
rect -1213 1320 -1212 2040
rect -492 1320 -491 2040
rect -1213 1319 -491 1320
rect -1632 1252 -1536 1268
rect -220 1268 -204 2092
rect -140 1268 -124 2092
rect 1192 2092 1288 2108
rect 199 2040 921 2041
rect 199 1320 200 2040
rect 920 1320 921 2040
rect 199 1319 921 1320
rect -220 1252 -124 1268
rect 1192 1268 1208 2092
rect 1272 1268 1288 2092
rect 2604 2092 2700 2108
rect 1611 2040 2333 2041
rect 1611 1320 1612 2040
rect 2332 1320 2333 2040
rect 1611 1319 2333 1320
rect 1192 1252 1288 1268
rect 2604 1268 2620 2092
rect 2684 1268 2700 2092
rect 4016 2092 4112 2108
rect 3023 2040 3745 2041
rect 3023 1320 3024 2040
rect 3744 1320 3745 2040
rect 3023 1319 3745 1320
rect 2604 1252 2700 1268
rect 4016 1268 4032 2092
rect 4096 1268 4112 2092
rect 5428 2092 5524 2108
rect 4435 2040 5157 2041
rect 4435 1320 4436 2040
rect 5156 1320 5157 2040
rect 4435 1319 5157 1320
rect 4016 1252 4112 1268
rect 5428 1268 5444 2092
rect 5508 1268 5524 2092
rect 6840 2092 6936 2108
rect 5847 2040 6569 2041
rect 5847 1320 5848 2040
rect 6568 1320 6569 2040
rect 5847 1319 6569 1320
rect 5428 1252 5524 1268
rect 6840 1268 6856 2092
rect 6920 1268 6936 2092
rect 8252 2092 8348 2108
rect 7259 2040 7981 2041
rect 7259 1320 7260 2040
rect 7980 1320 7981 2040
rect 7259 1319 7981 1320
rect 6840 1252 6936 1268
rect 8252 1268 8268 2092
rect 8332 1268 8348 2092
rect 9664 2092 9760 2108
rect 8671 2040 9393 2041
rect 8671 1320 8672 2040
rect 9392 1320 9393 2040
rect 8671 1319 9393 1320
rect 8252 1252 8348 1268
rect 9664 1268 9680 2092
rect 9744 1268 9760 2092
rect 11076 2092 11172 2108
rect 10083 2040 10805 2041
rect 10083 1320 10084 2040
rect 10804 1320 10805 2040
rect 10083 1319 10805 1320
rect 9664 1252 9760 1268
rect 11076 1268 11092 2092
rect 11156 1268 11172 2092
rect 12488 2092 12584 2108
rect 11495 2040 12217 2041
rect 11495 1320 11496 2040
rect 12216 1320 12217 2040
rect 11495 1319 12217 1320
rect 11076 1252 11172 1268
rect 12488 1268 12504 2092
rect 12568 1268 12584 2092
rect 13900 2092 13996 2108
rect 12907 2040 13629 2041
rect 12907 1320 12908 2040
rect 13628 1320 13629 2040
rect 12907 1319 13629 1320
rect 12488 1252 12584 1268
rect 13900 1268 13916 2092
rect 13980 1268 13996 2092
rect 15312 2092 15408 2108
rect 14319 2040 15041 2041
rect 14319 1320 14320 2040
rect 15040 1320 15041 2040
rect 14319 1319 15041 1320
rect 13900 1252 13996 1268
rect 15312 1268 15328 2092
rect 15392 1268 15408 2092
rect 16724 2092 16820 2108
rect 15731 2040 16453 2041
rect 15731 1320 15732 2040
rect 16452 1320 16453 2040
rect 15731 1319 16453 1320
rect 15312 1252 15408 1268
rect 16724 1268 16740 2092
rect 16804 1268 16820 2092
rect 18136 2092 18232 2108
rect 17143 2040 17865 2041
rect 17143 1320 17144 2040
rect 17864 1320 17865 2040
rect 17143 1319 17865 1320
rect 16724 1252 16820 1268
rect 18136 1268 18152 2092
rect 18216 1268 18232 2092
rect 19548 2092 19644 2108
rect 18555 2040 19277 2041
rect 18555 1320 18556 2040
rect 19276 1320 19277 2040
rect 18555 1319 19277 1320
rect 18136 1252 18232 1268
rect 19548 1268 19564 2092
rect 19628 1268 19644 2092
rect 20960 2092 21056 2108
rect 19967 2040 20689 2041
rect 19967 1320 19968 2040
rect 20688 1320 20689 2040
rect 19967 1319 20689 1320
rect 19548 1252 19644 1268
rect 20960 1268 20976 2092
rect 21040 1268 21056 2092
rect 22372 2092 22468 2108
rect 21379 2040 22101 2041
rect 21379 1320 21380 2040
rect 22100 1320 22101 2040
rect 21379 1319 22101 1320
rect 20960 1252 21056 1268
rect 22372 1268 22388 2092
rect 22452 1268 22468 2092
rect 23784 2092 23880 2108
rect 22791 2040 23513 2041
rect 22791 1320 22792 2040
rect 23512 1320 23513 2040
rect 22791 1319 23513 1320
rect 22372 1252 22468 1268
rect 23784 1268 23800 2092
rect 23864 1268 23880 2092
rect 23784 1252 23880 1268
rect -22812 972 -22716 988
rect -23805 920 -23083 921
rect -23805 200 -23804 920
rect -23084 200 -23083 920
rect -23805 199 -23083 200
rect -22812 148 -22796 972
rect -22732 148 -22716 972
rect -21400 972 -21304 988
rect -22393 920 -21671 921
rect -22393 200 -22392 920
rect -21672 200 -21671 920
rect -22393 199 -21671 200
rect -22812 132 -22716 148
rect -21400 148 -21384 972
rect -21320 148 -21304 972
rect -19988 972 -19892 988
rect -20981 920 -20259 921
rect -20981 200 -20980 920
rect -20260 200 -20259 920
rect -20981 199 -20259 200
rect -21400 132 -21304 148
rect -19988 148 -19972 972
rect -19908 148 -19892 972
rect -18576 972 -18480 988
rect -19569 920 -18847 921
rect -19569 200 -19568 920
rect -18848 200 -18847 920
rect -19569 199 -18847 200
rect -19988 132 -19892 148
rect -18576 148 -18560 972
rect -18496 148 -18480 972
rect -17164 972 -17068 988
rect -18157 920 -17435 921
rect -18157 200 -18156 920
rect -17436 200 -17435 920
rect -18157 199 -17435 200
rect -18576 132 -18480 148
rect -17164 148 -17148 972
rect -17084 148 -17068 972
rect -15752 972 -15656 988
rect -16745 920 -16023 921
rect -16745 200 -16744 920
rect -16024 200 -16023 920
rect -16745 199 -16023 200
rect -17164 132 -17068 148
rect -15752 148 -15736 972
rect -15672 148 -15656 972
rect -14340 972 -14244 988
rect -15333 920 -14611 921
rect -15333 200 -15332 920
rect -14612 200 -14611 920
rect -15333 199 -14611 200
rect -15752 132 -15656 148
rect -14340 148 -14324 972
rect -14260 148 -14244 972
rect -12928 972 -12832 988
rect -13921 920 -13199 921
rect -13921 200 -13920 920
rect -13200 200 -13199 920
rect -13921 199 -13199 200
rect -14340 132 -14244 148
rect -12928 148 -12912 972
rect -12848 148 -12832 972
rect -11516 972 -11420 988
rect -12509 920 -11787 921
rect -12509 200 -12508 920
rect -11788 200 -11787 920
rect -12509 199 -11787 200
rect -12928 132 -12832 148
rect -11516 148 -11500 972
rect -11436 148 -11420 972
rect -10104 972 -10008 988
rect -11097 920 -10375 921
rect -11097 200 -11096 920
rect -10376 200 -10375 920
rect -11097 199 -10375 200
rect -11516 132 -11420 148
rect -10104 148 -10088 972
rect -10024 148 -10008 972
rect -8692 972 -8596 988
rect -9685 920 -8963 921
rect -9685 200 -9684 920
rect -8964 200 -8963 920
rect -9685 199 -8963 200
rect -10104 132 -10008 148
rect -8692 148 -8676 972
rect -8612 148 -8596 972
rect -7280 972 -7184 988
rect -8273 920 -7551 921
rect -8273 200 -8272 920
rect -7552 200 -7551 920
rect -8273 199 -7551 200
rect -8692 132 -8596 148
rect -7280 148 -7264 972
rect -7200 148 -7184 972
rect -5868 972 -5772 988
rect -6861 920 -6139 921
rect -6861 200 -6860 920
rect -6140 200 -6139 920
rect -6861 199 -6139 200
rect -7280 132 -7184 148
rect -5868 148 -5852 972
rect -5788 148 -5772 972
rect -4456 972 -4360 988
rect -5449 920 -4727 921
rect -5449 200 -5448 920
rect -4728 200 -4727 920
rect -5449 199 -4727 200
rect -5868 132 -5772 148
rect -4456 148 -4440 972
rect -4376 148 -4360 972
rect -3044 972 -2948 988
rect -4037 920 -3315 921
rect -4037 200 -4036 920
rect -3316 200 -3315 920
rect -4037 199 -3315 200
rect -4456 132 -4360 148
rect -3044 148 -3028 972
rect -2964 148 -2948 972
rect -1632 972 -1536 988
rect -2625 920 -1903 921
rect -2625 200 -2624 920
rect -1904 200 -1903 920
rect -2625 199 -1903 200
rect -3044 132 -2948 148
rect -1632 148 -1616 972
rect -1552 148 -1536 972
rect -220 972 -124 988
rect -1213 920 -491 921
rect -1213 200 -1212 920
rect -492 200 -491 920
rect -1213 199 -491 200
rect -1632 132 -1536 148
rect -220 148 -204 972
rect -140 148 -124 972
rect 1192 972 1288 988
rect 199 920 921 921
rect 199 200 200 920
rect 920 200 921 920
rect 199 199 921 200
rect -220 132 -124 148
rect 1192 148 1208 972
rect 1272 148 1288 972
rect 2604 972 2700 988
rect 1611 920 2333 921
rect 1611 200 1612 920
rect 2332 200 2333 920
rect 1611 199 2333 200
rect 1192 132 1288 148
rect 2604 148 2620 972
rect 2684 148 2700 972
rect 4016 972 4112 988
rect 3023 920 3745 921
rect 3023 200 3024 920
rect 3744 200 3745 920
rect 3023 199 3745 200
rect 2604 132 2700 148
rect 4016 148 4032 972
rect 4096 148 4112 972
rect 5428 972 5524 988
rect 4435 920 5157 921
rect 4435 200 4436 920
rect 5156 200 5157 920
rect 4435 199 5157 200
rect 4016 132 4112 148
rect 5428 148 5444 972
rect 5508 148 5524 972
rect 6840 972 6936 988
rect 5847 920 6569 921
rect 5847 200 5848 920
rect 6568 200 6569 920
rect 5847 199 6569 200
rect 5428 132 5524 148
rect 6840 148 6856 972
rect 6920 148 6936 972
rect 8252 972 8348 988
rect 7259 920 7981 921
rect 7259 200 7260 920
rect 7980 200 7981 920
rect 7259 199 7981 200
rect 6840 132 6936 148
rect 8252 148 8268 972
rect 8332 148 8348 972
rect 9664 972 9760 988
rect 8671 920 9393 921
rect 8671 200 8672 920
rect 9392 200 9393 920
rect 8671 199 9393 200
rect 8252 132 8348 148
rect 9664 148 9680 972
rect 9744 148 9760 972
rect 11076 972 11172 988
rect 10083 920 10805 921
rect 10083 200 10084 920
rect 10804 200 10805 920
rect 10083 199 10805 200
rect 9664 132 9760 148
rect 11076 148 11092 972
rect 11156 148 11172 972
rect 12488 972 12584 988
rect 11495 920 12217 921
rect 11495 200 11496 920
rect 12216 200 12217 920
rect 11495 199 12217 200
rect 11076 132 11172 148
rect 12488 148 12504 972
rect 12568 148 12584 972
rect 13900 972 13996 988
rect 12907 920 13629 921
rect 12907 200 12908 920
rect 13628 200 13629 920
rect 12907 199 13629 200
rect 12488 132 12584 148
rect 13900 148 13916 972
rect 13980 148 13996 972
rect 15312 972 15408 988
rect 14319 920 15041 921
rect 14319 200 14320 920
rect 15040 200 15041 920
rect 14319 199 15041 200
rect 13900 132 13996 148
rect 15312 148 15328 972
rect 15392 148 15408 972
rect 16724 972 16820 988
rect 15731 920 16453 921
rect 15731 200 15732 920
rect 16452 200 16453 920
rect 15731 199 16453 200
rect 15312 132 15408 148
rect 16724 148 16740 972
rect 16804 148 16820 972
rect 18136 972 18232 988
rect 17143 920 17865 921
rect 17143 200 17144 920
rect 17864 200 17865 920
rect 17143 199 17865 200
rect 16724 132 16820 148
rect 18136 148 18152 972
rect 18216 148 18232 972
rect 19548 972 19644 988
rect 18555 920 19277 921
rect 18555 200 18556 920
rect 19276 200 19277 920
rect 18555 199 19277 200
rect 18136 132 18232 148
rect 19548 148 19564 972
rect 19628 148 19644 972
rect 20960 972 21056 988
rect 19967 920 20689 921
rect 19967 200 19968 920
rect 20688 200 20689 920
rect 19967 199 20689 200
rect 19548 132 19644 148
rect 20960 148 20976 972
rect 21040 148 21056 972
rect 22372 972 22468 988
rect 21379 920 22101 921
rect 21379 200 21380 920
rect 22100 200 22101 920
rect 21379 199 22101 200
rect 20960 132 21056 148
rect 22372 148 22388 972
rect 22452 148 22468 972
rect 23784 972 23880 988
rect 22791 920 23513 921
rect 22791 200 22792 920
rect 23512 200 23513 920
rect 22791 199 23513 200
rect 22372 132 22468 148
rect 23784 148 23800 972
rect 23864 148 23880 972
rect 23784 132 23880 148
rect -22812 -148 -22716 -132
rect -23805 -200 -23083 -199
rect -23805 -920 -23804 -200
rect -23084 -920 -23083 -200
rect -23805 -921 -23083 -920
rect -22812 -972 -22796 -148
rect -22732 -972 -22716 -148
rect -21400 -148 -21304 -132
rect -22393 -200 -21671 -199
rect -22393 -920 -22392 -200
rect -21672 -920 -21671 -200
rect -22393 -921 -21671 -920
rect -22812 -988 -22716 -972
rect -21400 -972 -21384 -148
rect -21320 -972 -21304 -148
rect -19988 -148 -19892 -132
rect -20981 -200 -20259 -199
rect -20981 -920 -20980 -200
rect -20260 -920 -20259 -200
rect -20981 -921 -20259 -920
rect -21400 -988 -21304 -972
rect -19988 -972 -19972 -148
rect -19908 -972 -19892 -148
rect -18576 -148 -18480 -132
rect -19569 -200 -18847 -199
rect -19569 -920 -19568 -200
rect -18848 -920 -18847 -200
rect -19569 -921 -18847 -920
rect -19988 -988 -19892 -972
rect -18576 -972 -18560 -148
rect -18496 -972 -18480 -148
rect -17164 -148 -17068 -132
rect -18157 -200 -17435 -199
rect -18157 -920 -18156 -200
rect -17436 -920 -17435 -200
rect -18157 -921 -17435 -920
rect -18576 -988 -18480 -972
rect -17164 -972 -17148 -148
rect -17084 -972 -17068 -148
rect -15752 -148 -15656 -132
rect -16745 -200 -16023 -199
rect -16745 -920 -16744 -200
rect -16024 -920 -16023 -200
rect -16745 -921 -16023 -920
rect -17164 -988 -17068 -972
rect -15752 -972 -15736 -148
rect -15672 -972 -15656 -148
rect -14340 -148 -14244 -132
rect -15333 -200 -14611 -199
rect -15333 -920 -15332 -200
rect -14612 -920 -14611 -200
rect -15333 -921 -14611 -920
rect -15752 -988 -15656 -972
rect -14340 -972 -14324 -148
rect -14260 -972 -14244 -148
rect -12928 -148 -12832 -132
rect -13921 -200 -13199 -199
rect -13921 -920 -13920 -200
rect -13200 -920 -13199 -200
rect -13921 -921 -13199 -920
rect -14340 -988 -14244 -972
rect -12928 -972 -12912 -148
rect -12848 -972 -12832 -148
rect -11516 -148 -11420 -132
rect -12509 -200 -11787 -199
rect -12509 -920 -12508 -200
rect -11788 -920 -11787 -200
rect -12509 -921 -11787 -920
rect -12928 -988 -12832 -972
rect -11516 -972 -11500 -148
rect -11436 -972 -11420 -148
rect -10104 -148 -10008 -132
rect -11097 -200 -10375 -199
rect -11097 -920 -11096 -200
rect -10376 -920 -10375 -200
rect -11097 -921 -10375 -920
rect -11516 -988 -11420 -972
rect -10104 -972 -10088 -148
rect -10024 -972 -10008 -148
rect -8692 -148 -8596 -132
rect -9685 -200 -8963 -199
rect -9685 -920 -9684 -200
rect -8964 -920 -8963 -200
rect -9685 -921 -8963 -920
rect -10104 -988 -10008 -972
rect -8692 -972 -8676 -148
rect -8612 -972 -8596 -148
rect -7280 -148 -7184 -132
rect -8273 -200 -7551 -199
rect -8273 -920 -8272 -200
rect -7552 -920 -7551 -200
rect -8273 -921 -7551 -920
rect -8692 -988 -8596 -972
rect -7280 -972 -7264 -148
rect -7200 -972 -7184 -148
rect -5868 -148 -5772 -132
rect -6861 -200 -6139 -199
rect -6861 -920 -6860 -200
rect -6140 -920 -6139 -200
rect -6861 -921 -6139 -920
rect -7280 -988 -7184 -972
rect -5868 -972 -5852 -148
rect -5788 -972 -5772 -148
rect -4456 -148 -4360 -132
rect -5449 -200 -4727 -199
rect -5449 -920 -5448 -200
rect -4728 -920 -4727 -200
rect -5449 -921 -4727 -920
rect -5868 -988 -5772 -972
rect -4456 -972 -4440 -148
rect -4376 -972 -4360 -148
rect -3044 -148 -2948 -132
rect -4037 -200 -3315 -199
rect -4037 -920 -4036 -200
rect -3316 -920 -3315 -200
rect -4037 -921 -3315 -920
rect -4456 -988 -4360 -972
rect -3044 -972 -3028 -148
rect -2964 -972 -2948 -148
rect -1632 -148 -1536 -132
rect -2625 -200 -1903 -199
rect -2625 -920 -2624 -200
rect -1904 -920 -1903 -200
rect -2625 -921 -1903 -920
rect -3044 -988 -2948 -972
rect -1632 -972 -1616 -148
rect -1552 -972 -1536 -148
rect -220 -148 -124 -132
rect -1213 -200 -491 -199
rect -1213 -920 -1212 -200
rect -492 -920 -491 -200
rect -1213 -921 -491 -920
rect -1632 -988 -1536 -972
rect -220 -972 -204 -148
rect -140 -972 -124 -148
rect 1192 -148 1288 -132
rect 199 -200 921 -199
rect 199 -920 200 -200
rect 920 -920 921 -200
rect 199 -921 921 -920
rect -220 -988 -124 -972
rect 1192 -972 1208 -148
rect 1272 -972 1288 -148
rect 2604 -148 2700 -132
rect 1611 -200 2333 -199
rect 1611 -920 1612 -200
rect 2332 -920 2333 -200
rect 1611 -921 2333 -920
rect 1192 -988 1288 -972
rect 2604 -972 2620 -148
rect 2684 -972 2700 -148
rect 4016 -148 4112 -132
rect 3023 -200 3745 -199
rect 3023 -920 3024 -200
rect 3744 -920 3745 -200
rect 3023 -921 3745 -920
rect 2604 -988 2700 -972
rect 4016 -972 4032 -148
rect 4096 -972 4112 -148
rect 5428 -148 5524 -132
rect 4435 -200 5157 -199
rect 4435 -920 4436 -200
rect 5156 -920 5157 -200
rect 4435 -921 5157 -920
rect 4016 -988 4112 -972
rect 5428 -972 5444 -148
rect 5508 -972 5524 -148
rect 6840 -148 6936 -132
rect 5847 -200 6569 -199
rect 5847 -920 5848 -200
rect 6568 -920 6569 -200
rect 5847 -921 6569 -920
rect 5428 -988 5524 -972
rect 6840 -972 6856 -148
rect 6920 -972 6936 -148
rect 8252 -148 8348 -132
rect 7259 -200 7981 -199
rect 7259 -920 7260 -200
rect 7980 -920 7981 -200
rect 7259 -921 7981 -920
rect 6840 -988 6936 -972
rect 8252 -972 8268 -148
rect 8332 -972 8348 -148
rect 9664 -148 9760 -132
rect 8671 -200 9393 -199
rect 8671 -920 8672 -200
rect 9392 -920 9393 -200
rect 8671 -921 9393 -920
rect 8252 -988 8348 -972
rect 9664 -972 9680 -148
rect 9744 -972 9760 -148
rect 11076 -148 11172 -132
rect 10083 -200 10805 -199
rect 10083 -920 10084 -200
rect 10804 -920 10805 -200
rect 10083 -921 10805 -920
rect 9664 -988 9760 -972
rect 11076 -972 11092 -148
rect 11156 -972 11172 -148
rect 12488 -148 12584 -132
rect 11495 -200 12217 -199
rect 11495 -920 11496 -200
rect 12216 -920 12217 -200
rect 11495 -921 12217 -920
rect 11076 -988 11172 -972
rect 12488 -972 12504 -148
rect 12568 -972 12584 -148
rect 13900 -148 13996 -132
rect 12907 -200 13629 -199
rect 12907 -920 12908 -200
rect 13628 -920 13629 -200
rect 12907 -921 13629 -920
rect 12488 -988 12584 -972
rect 13900 -972 13916 -148
rect 13980 -972 13996 -148
rect 15312 -148 15408 -132
rect 14319 -200 15041 -199
rect 14319 -920 14320 -200
rect 15040 -920 15041 -200
rect 14319 -921 15041 -920
rect 13900 -988 13996 -972
rect 15312 -972 15328 -148
rect 15392 -972 15408 -148
rect 16724 -148 16820 -132
rect 15731 -200 16453 -199
rect 15731 -920 15732 -200
rect 16452 -920 16453 -200
rect 15731 -921 16453 -920
rect 15312 -988 15408 -972
rect 16724 -972 16740 -148
rect 16804 -972 16820 -148
rect 18136 -148 18232 -132
rect 17143 -200 17865 -199
rect 17143 -920 17144 -200
rect 17864 -920 17865 -200
rect 17143 -921 17865 -920
rect 16724 -988 16820 -972
rect 18136 -972 18152 -148
rect 18216 -972 18232 -148
rect 19548 -148 19644 -132
rect 18555 -200 19277 -199
rect 18555 -920 18556 -200
rect 19276 -920 19277 -200
rect 18555 -921 19277 -920
rect 18136 -988 18232 -972
rect 19548 -972 19564 -148
rect 19628 -972 19644 -148
rect 20960 -148 21056 -132
rect 19967 -200 20689 -199
rect 19967 -920 19968 -200
rect 20688 -920 20689 -200
rect 19967 -921 20689 -920
rect 19548 -988 19644 -972
rect 20960 -972 20976 -148
rect 21040 -972 21056 -148
rect 22372 -148 22468 -132
rect 21379 -200 22101 -199
rect 21379 -920 21380 -200
rect 22100 -920 22101 -200
rect 21379 -921 22101 -920
rect 20960 -988 21056 -972
rect 22372 -972 22388 -148
rect 22452 -972 22468 -148
rect 23784 -148 23880 -132
rect 22791 -200 23513 -199
rect 22791 -920 22792 -200
rect 23512 -920 23513 -200
rect 22791 -921 23513 -920
rect 22372 -988 22468 -972
rect 23784 -972 23800 -148
rect 23864 -972 23880 -148
rect 23784 -988 23880 -972
rect -22812 -1268 -22716 -1252
rect -23805 -1320 -23083 -1319
rect -23805 -2040 -23804 -1320
rect -23084 -2040 -23083 -1320
rect -23805 -2041 -23083 -2040
rect -22812 -2092 -22796 -1268
rect -22732 -2092 -22716 -1268
rect -21400 -1268 -21304 -1252
rect -22393 -1320 -21671 -1319
rect -22393 -2040 -22392 -1320
rect -21672 -2040 -21671 -1320
rect -22393 -2041 -21671 -2040
rect -22812 -2108 -22716 -2092
rect -21400 -2092 -21384 -1268
rect -21320 -2092 -21304 -1268
rect -19988 -1268 -19892 -1252
rect -20981 -1320 -20259 -1319
rect -20981 -2040 -20980 -1320
rect -20260 -2040 -20259 -1320
rect -20981 -2041 -20259 -2040
rect -21400 -2108 -21304 -2092
rect -19988 -2092 -19972 -1268
rect -19908 -2092 -19892 -1268
rect -18576 -1268 -18480 -1252
rect -19569 -1320 -18847 -1319
rect -19569 -2040 -19568 -1320
rect -18848 -2040 -18847 -1320
rect -19569 -2041 -18847 -2040
rect -19988 -2108 -19892 -2092
rect -18576 -2092 -18560 -1268
rect -18496 -2092 -18480 -1268
rect -17164 -1268 -17068 -1252
rect -18157 -1320 -17435 -1319
rect -18157 -2040 -18156 -1320
rect -17436 -2040 -17435 -1320
rect -18157 -2041 -17435 -2040
rect -18576 -2108 -18480 -2092
rect -17164 -2092 -17148 -1268
rect -17084 -2092 -17068 -1268
rect -15752 -1268 -15656 -1252
rect -16745 -1320 -16023 -1319
rect -16745 -2040 -16744 -1320
rect -16024 -2040 -16023 -1320
rect -16745 -2041 -16023 -2040
rect -17164 -2108 -17068 -2092
rect -15752 -2092 -15736 -1268
rect -15672 -2092 -15656 -1268
rect -14340 -1268 -14244 -1252
rect -15333 -1320 -14611 -1319
rect -15333 -2040 -15332 -1320
rect -14612 -2040 -14611 -1320
rect -15333 -2041 -14611 -2040
rect -15752 -2108 -15656 -2092
rect -14340 -2092 -14324 -1268
rect -14260 -2092 -14244 -1268
rect -12928 -1268 -12832 -1252
rect -13921 -1320 -13199 -1319
rect -13921 -2040 -13920 -1320
rect -13200 -2040 -13199 -1320
rect -13921 -2041 -13199 -2040
rect -14340 -2108 -14244 -2092
rect -12928 -2092 -12912 -1268
rect -12848 -2092 -12832 -1268
rect -11516 -1268 -11420 -1252
rect -12509 -1320 -11787 -1319
rect -12509 -2040 -12508 -1320
rect -11788 -2040 -11787 -1320
rect -12509 -2041 -11787 -2040
rect -12928 -2108 -12832 -2092
rect -11516 -2092 -11500 -1268
rect -11436 -2092 -11420 -1268
rect -10104 -1268 -10008 -1252
rect -11097 -1320 -10375 -1319
rect -11097 -2040 -11096 -1320
rect -10376 -2040 -10375 -1320
rect -11097 -2041 -10375 -2040
rect -11516 -2108 -11420 -2092
rect -10104 -2092 -10088 -1268
rect -10024 -2092 -10008 -1268
rect -8692 -1268 -8596 -1252
rect -9685 -1320 -8963 -1319
rect -9685 -2040 -9684 -1320
rect -8964 -2040 -8963 -1320
rect -9685 -2041 -8963 -2040
rect -10104 -2108 -10008 -2092
rect -8692 -2092 -8676 -1268
rect -8612 -2092 -8596 -1268
rect -7280 -1268 -7184 -1252
rect -8273 -1320 -7551 -1319
rect -8273 -2040 -8272 -1320
rect -7552 -2040 -7551 -1320
rect -8273 -2041 -7551 -2040
rect -8692 -2108 -8596 -2092
rect -7280 -2092 -7264 -1268
rect -7200 -2092 -7184 -1268
rect -5868 -1268 -5772 -1252
rect -6861 -1320 -6139 -1319
rect -6861 -2040 -6860 -1320
rect -6140 -2040 -6139 -1320
rect -6861 -2041 -6139 -2040
rect -7280 -2108 -7184 -2092
rect -5868 -2092 -5852 -1268
rect -5788 -2092 -5772 -1268
rect -4456 -1268 -4360 -1252
rect -5449 -1320 -4727 -1319
rect -5449 -2040 -5448 -1320
rect -4728 -2040 -4727 -1320
rect -5449 -2041 -4727 -2040
rect -5868 -2108 -5772 -2092
rect -4456 -2092 -4440 -1268
rect -4376 -2092 -4360 -1268
rect -3044 -1268 -2948 -1252
rect -4037 -1320 -3315 -1319
rect -4037 -2040 -4036 -1320
rect -3316 -2040 -3315 -1320
rect -4037 -2041 -3315 -2040
rect -4456 -2108 -4360 -2092
rect -3044 -2092 -3028 -1268
rect -2964 -2092 -2948 -1268
rect -1632 -1268 -1536 -1252
rect -2625 -1320 -1903 -1319
rect -2625 -2040 -2624 -1320
rect -1904 -2040 -1903 -1320
rect -2625 -2041 -1903 -2040
rect -3044 -2108 -2948 -2092
rect -1632 -2092 -1616 -1268
rect -1552 -2092 -1536 -1268
rect -220 -1268 -124 -1252
rect -1213 -1320 -491 -1319
rect -1213 -2040 -1212 -1320
rect -492 -2040 -491 -1320
rect -1213 -2041 -491 -2040
rect -1632 -2108 -1536 -2092
rect -220 -2092 -204 -1268
rect -140 -2092 -124 -1268
rect 1192 -1268 1288 -1252
rect 199 -1320 921 -1319
rect 199 -2040 200 -1320
rect 920 -2040 921 -1320
rect 199 -2041 921 -2040
rect -220 -2108 -124 -2092
rect 1192 -2092 1208 -1268
rect 1272 -2092 1288 -1268
rect 2604 -1268 2700 -1252
rect 1611 -1320 2333 -1319
rect 1611 -2040 1612 -1320
rect 2332 -2040 2333 -1320
rect 1611 -2041 2333 -2040
rect 1192 -2108 1288 -2092
rect 2604 -2092 2620 -1268
rect 2684 -2092 2700 -1268
rect 4016 -1268 4112 -1252
rect 3023 -1320 3745 -1319
rect 3023 -2040 3024 -1320
rect 3744 -2040 3745 -1320
rect 3023 -2041 3745 -2040
rect 2604 -2108 2700 -2092
rect 4016 -2092 4032 -1268
rect 4096 -2092 4112 -1268
rect 5428 -1268 5524 -1252
rect 4435 -1320 5157 -1319
rect 4435 -2040 4436 -1320
rect 5156 -2040 5157 -1320
rect 4435 -2041 5157 -2040
rect 4016 -2108 4112 -2092
rect 5428 -2092 5444 -1268
rect 5508 -2092 5524 -1268
rect 6840 -1268 6936 -1252
rect 5847 -1320 6569 -1319
rect 5847 -2040 5848 -1320
rect 6568 -2040 6569 -1320
rect 5847 -2041 6569 -2040
rect 5428 -2108 5524 -2092
rect 6840 -2092 6856 -1268
rect 6920 -2092 6936 -1268
rect 8252 -1268 8348 -1252
rect 7259 -1320 7981 -1319
rect 7259 -2040 7260 -1320
rect 7980 -2040 7981 -1320
rect 7259 -2041 7981 -2040
rect 6840 -2108 6936 -2092
rect 8252 -2092 8268 -1268
rect 8332 -2092 8348 -1268
rect 9664 -1268 9760 -1252
rect 8671 -1320 9393 -1319
rect 8671 -2040 8672 -1320
rect 9392 -2040 9393 -1320
rect 8671 -2041 9393 -2040
rect 8252 -2108 8348 -2092
rect 9664 -2092 9680 -1268
rect 9744 -2092 9760 -1268
rect 11076 -1268 11172 -1252
rect 10083 -1320 10805 -1319
rect 10083 -2040 10084 -1320
rect 10804 -2040 10805 -1320
rect 10083 -2041 10805 -2040
rect 9664 -2108 9760 -2092
rect 11076 -2092 11092 -1268
rect 11156 -2092 11172 -1268
rect 12488 -1268 12584 -1252
rect 11495 -1320 12217 -1319
rect 11495 -2040 11496 -1320
rect 12216 -2040 12217 -1320
rect 11495 -2041 12217 -2040
rect 11076 -2108 11172 -2092
rect 12488 -2092 12504 -1268
rect 12568 -2092 12584 -1268
rect 13900 -1268 13996 -1252
rect 12907 -1320 13629 -1319
rect 12907 -2040 12908 -1320
rect 13628 -2040 13629 -1320
rect 12907 -2041 13629 -2040
rect 12488 -2108 12584 -2092
rect 13900 -2092 13916 -1268
rect 13980 -2092 13996 -1268
rect 15312 -1268 15408 -1252
rect 14319 -1320 15041 -1319
rect 14319 -2040 14320 -1320
rect 15040 -2040 15041 -1320
rect 14319 -2041 15041 -2040
rect 13900 -2108 13996 -2092
rect 15312 -2092 15328 -1268
rect 15392 -2092 15408 -1268
rect 16724 -1268 16820 -1252
rect 15731 -1320 16453 -1319
rect 15731 -2040 15732 -1320
rect 16452 -2040 16453 -1320
rect 15731 -2041 16453 -2040
rect 15312 -2108 15408 -2092
rect 16724 -2092 16740 -1268
rect 16804 -2092 16820 -1268
rect 18136 -1268 18232 -1252
rect 17143 -1320 17865 -1319
rect 17143 -2040 17144 -1320
rect 17864 -2040 17865 -1320
rect 17143 -2041 17865 -2040
rect 16724 -2108 16820 -2092
rect 18136 -2092 18152 -1268
rect 18216 -2092 18232 -1268
rect 19548 -1268 19644 -1252
rect 18555 -1320 19277 -1319
rect 18555 -2040 18556 -1320
rect 19276 -2040 19277 -1320
rect 18555 -2041 19277 -2040
rect 18136 -2108 18232 -2092
rect 19548 -2092 19564 -1268
rect 19628 -2092 19644 -1268
rect 20960 -1268 21056 -1252
rect 19967 -1320 20689 -1319
rect 19967 -2040 19968 -1320
rect 20688 -2040 20689 -1320
rect 19967 -2041 20689 -2040
rect 19548 -2108 19644 -2092
rect 20960 -2092 20976 -1268
rect 21040 -2092 21056 -1268
rect 22372 -1268 22468 -1252
rect 21379 -1320 22101 -1319
rect 21379 -2040 21380 -1320
rect 22100 -2040 22101 -1320
rect 21379 -2041 22101 -2040
rect 20960 -2108 21056 -2092
rect 22372 -2092 22388 -1268
rect 22452 -2092 22468 -1268
rect 23784 -1268 23880 -1252
rect 22791 -1320 23513 -1319
rect 22791 -2040 22792 -1320
rect 23512 -2040 23513 -1320
rect 22791 -2041 23513 -2040
rect 22372 -2108 22468 -2092
rect 23784 -2092 23800 -1268
rect 23864 -2092 23880 -1268
rect 23784 -2108 23880 -2092
rect -22812 -2388 -22716 -2372
rect -23805 -2440 -23083 -2439
rect -23805 -3160 -23804 -2440
rect -23084 -3160 -23083 -2440
rect -23805 -3161 -23083 -3160
rect -22812 -3212 -22796 -2388
rect -22732 -3212 -22716 -2388
rect -21400 -2388 -21304 -2372
rect -22393 -2440 -21671 -2439
rect -22393 -3160 -22392 -2440
rect -21672 -3160 -21671 -2440
rect -22393 -3161 -21671 -3160
rect -22812 -3228 -22716 -3212
rect -21400 -3212 -21384 -2388
rect -21320 -3212 -21304 -2388
rect -19988 -2388 -19892 -2372
rect -20981 -2440 -20259 -2439
rect -20981 -3160 -20980 -2440
rect -20260 -3160 -20259 -2440
rect -20981 -3161 -20259 -3160
rect -21400 -3228 -21304 -3212
rect -19988 -3212 -19972 -2388
rect -19908 -3212 -19892 -2388
rect -18576 -2388 -18480 -2372
rect -19569 -2440 -18847 -2439
rect -19569 -3160 -19568 -2440
rect -18848 -3160 -18847 -2440
rect -19569 -3161 -18847 -3160
rect -19988 -3228 -19892 -3212
rect -18576 -3212 -18560 -2388
rect -18496 -3212 -18480 -2388
rect -17164 -2388 -17068 -2372
rect -18157 -2440 -17435 -2439
rect -18157 -3160 -18156 -2440
rect -17436 -3160 -17435 -2440
rect -18157 -3161 -17435 -3160
rect -18576 -3228 -18480 -3212
rect -17164 -3212 -17148 -2388
rect -17084 -3212 -17068 -2388
rect -15752 -2388 -15656 -2372
rect -16745 -2440 -16023 -2439
rect -16745 -3160 -16744 -2440
rect -16024 -3160 -16023 -2440
rect -16745 -3161 -16023 -3160
rect -17164 -3228 -17068 -3212
rect -15752 -3212 -15736 -2388
rect -15672 -3212 -15656 -2388
rect -14340 -2388 -14244 -2372
rect -15333 -2440 -14611 -2439
rect -15333 -3160 -15332 -2440
rect -14612 -3160 -14611 -2440
rect -15333 -3161 -14611 -3160
rect -15752 -3228 -15656 -3212
rect -14340 -3212 -14324 -2388
rect -14260 -3212 -14244 -2388
rect -12928 -2388 -12832 -2372
rect -13921 -2440 -13199 -2439
rect -13921 -3160 -13920 -2440
rect -13200 -3160 -13199 -2440
rect -13921 -3161 -13199 -3160
rect -14340 -3228 -14244 -3212
rect -12928 -3212 -12912 -2388
rect -12848 -3212 -12832 -2388
rect -11516 -2388 -11420 -2372
rect -12509 -2440 -11787 -2439
rect -12509 -3160 -12508 -2440
rect -11788 -3160 -11787 -2440
rect -12509 -3161 -11787 -3160
rect -12928 -3228 -12832 -3212
rect -11516 -3212 -11500 -2388
rect -11436 -3212 -11420 -2388
rect -10104 -2388 -10008 -2372
rect -11097 -2440 -10375 -2439
rect -11097 -3160 -11096 -2440
rect -10376 -3160 -10375 -2440
rect -11097 -3161 -10375 -3160
rect -11516 -3228 -11420 -3212
rect -10104 -3212 -10088 -2388
rect -10024 -3212 -10008 -2388
rect -8692 -2388 -8596 -2372
rect -9685 -2440 -8963 -2439
rect -9685 -3160 -9684 -2440
rect -8964 -3160 -8963 -2440
rect -9685 -3161 -8963 -3160
rect -10104 -3228 -10008 -3212
rect -8692 -3212 -8676 -2388
rect -8612 -3212 -8596 -2388
rect -7280 -2388 -7184 -2372
rect -8273 -2440 -7551 -2439
rect -8273 -3160 -8272 -2440
rect -7552 -3160 -7551 -2440
rect -8273 -3161 -7551 -3160
rect -8692 -3228 -8596 -3212
rect -7280 -3212 -7264 -2388
rect -7200 -3212 -7184 -2388
rect -5868 -2388 -5772 -2372
rect -6861 -2440 -6139 -2439
rect -6861 -3160 -6860 -2440
rect -6140 -3160 -6139 -2440
rect -6861 -3161 -6139 -3160
rect -7280 -3228 -7184 -3212
rect -5868 -3212 -5852 -2388
rect -5788 -3212 -5772 -2388
rect -4456 -2388 -4360 -2372
rect -5449 -2440 -4727 -2439
rect -5449 -3160 -5448 -2440
rect -4728 -3160 -4727 -2440
rect -5449 -3161 -4727 -3160
rect -5868 -3228 -5772 -3212
rect -4456 -3212 -4440 -2388
rect -4376 -3212 -4360 -2388
rect -3044 -2388 -2948 -2372
rect -4037 -2440 -3315 -2439
rect -4037 -3160 -4036 -2440
rect -3316 -3160 -3315 -2440
rect -4037 -3161 -3315 -3160
rect -4456 -3228 -4360 -3212
rect -3044 -3212 -3028 -2388
rect -2964 -3212 -2948 -2388
rect -1632 -2388 -1536 -2372
rect -2625 -2440 -1903 -2439
rect -2625 -3160 -2624 -2440
rect -1904 -3160 -1903 -2440
rect -2625 -3161 -1903 -3160
rect -3044 -3228 -2948 -3212
rect -1632 -3212 -1616 -2388
rect -1552 -3212 -1536 -2388
rect -220 -2388 -124 -2372
rect -1213 -2440 -491 -2439
rect -1213 -3160 -1212 -2440
rect -492 -3160 -491 -2440
rect -1213 -3161 -491 -3160
rect -1632 -3228 -1536 -3212
rect -220 -3212 -204 -2388
rect -140 -3212 -124 -2388
rect 1192 -2388 1288 -2372
rect 199 -2440 921 -2439
rect 199 -3160 200 -2440
rect 920 -3160 921 -2440
rect 199 -3161 921 -3160
rect -220 -3228 -124 -3212
rect 1192 -3212 1208 -2388
rect 1272 -3212 1288 -2388
rect 2604 -2388 2700 -2372
rect 1611 -2440 2333 -2439
rect 1611 -3160 1612 -2440
rect 2332 -3160 2333 -2440
rect 1611 -3161 2333 -3160
rect 1192 -3228 1288 -3212
rect 2604 -3212 2620 -2388
rect 2684 -3212 2700 -2388
rect 4016 -2388 4112 -2372
rect 3023 -2440 3745 -2439
rect 3023 -3160 3024 -2440
rect 3744 -3160 3745 -2440
rect 3023 -3161 3745 -3160
rect 2604 -3228 2700 -3212
rect 4016 -3212 4032 -2388
rect 4096 -3212 4112 -2388
rect 5428 -2388 5524 -2372
rect 4435 -2440 5157 -2439
rect 4435 -3160 4436 -2440
rect 5156 -3160 5157 -2440
rect 4435 -3161 5157 -3160
rect 4016 -3228 4112 -3212
rect 5428 -3212 5444 -2388
rect 5508 -3212 5524 -2388
rect 6840 -2388 6936 -2372
rect 5847 -2440 6569 -2439
rect 5847 -3160 5848 -2440
rect 6568 -3160 6569 -2440
rect 5847 -3161 6569 -3160
rect 5428 -3228 5524 -3212
rect 6840 -3212 6856 -2388
rect 6920 -3212 6936 -2388
rect 8252 -2388 8348 -2372
rect 7259 -2440 7981 -2439
rect 7259 -3160 7260 -2440
rect 7980 -3160 7981 -2440
rect 7259 -3161 7981 -3160
rect 6840 -3228 6936 -3212
rect 8252 -3212 8268 -2388
rect 8332 -3212 8348 -2388
rect 9664 -2388 9760 -2372
rect 8671 -2440 9393 -2439
rect 8671 -3160 8672 -2440
rect 9392 -3160 9393 -2440
rect 8671 -3161 9393 -3160
rect 8252 -3228 8348 -3212
rect 9664 -3212 9680 -2388
rect 9744 -3212 9760 -2388
rect 11076 -2388 11172 -2372
rect 10083 -2440 10805 -2439
rect 10083 -3160 10084 -2440
rect 10804 -3160 10805 -2440
rect 10083 -3161 10805 -3160
rect 9664 -3228 9760 -3212
rect 11076 -3212 11092 -2388
rect 11156 -3212 11172 -2388
rect 12488 -2388 12584 -2372
rect 11495 -2440 12217 -2439
rect 11495 -3160 11496 -2440
rect 12216 -3160 12217 -2440
rect 11495 -3161 12217 -3160
rect 11076 -3228 11172 -3212
rect 12488 -3212 12504 -2388
rect 12568 -3212 12584 -2388
rect 13900 -2388 13996 -2372
rect 12907 -2440 13629 -2439
rect 12907 -3160 12908 -2440
rect 13628 -3160 13629 -2440
rect 12907 -3161 13629 -3160
rect 12488 -3228 12584 -3212
rect 13900 -3212 13916 -2388
rect 13980 -3212 13996 -2388
rect 15312 -2388 15408 -2372
rect 14319 -2440 15041 -2439
rect 14319 -3160 14320 -2440
rect 15040 -3160 15041 -2440
rect 14319 -3161 15041 -3160
rect 13900 -3228 13996 -3212
rect 15312 -3212 15328 -2388
rect 15392 -3212 15408 -2388
rect 16724 -2388 16820 -2372
rect 15731 -2440 16453 -2439
rect 15731 -3160 15732 -2440
rect 16452 -3160 16453 -2440
rect 15731 -3161 16453 -3160
rect 15312 -3228 15408 -3212
rect 16724 -3212 16740 -2388
rect 16804 -3212 16820 -2388
rect 18136 -2388 18232 -2372
rect 17143 -2440 17865 -2439
rect 17143 -3160 17144 -2440
rect 17864 -3160 17865 -2440
rect 17143 -3161 17865 -3160
rect 16724 -3228 16820 -3212
rect 18136 -3212 18152 -2388
rect 18216 -3212 18232 -2388
rect 19548 -2388 19644 -2372
rect 18555 -2440 19277 -2439
rect 18555 -3160 18556 -2440
rect 19276 -3160 19277 -2440
rect 18555 -3161 19277 -3160
rect 18136 -3228 18232 -3212
rect 19548 -3212 19564 -2388
rect 19628 -3212 19644 -2388
rect 20960 -2388 21056 -2372
rect 19967 -2440 20689 -2439
rect 19967 -3160 19968 -2440
rect 20688 -3160 20689 -2440
rect 19967 -3161 20689 -3160
rect 19548 -3228 19644 -3212
rect 20960 -3212 20976 -2388
rect 21040 -3212 21056 -2388
rect 22372 -2388 22468 -2372
rect 21379 -2440 22101 -2439
rect 21379 -3160 21380 -2440
rect 22100 -3160 22101 -2440
rect 21379 -3161 22101 -3160
rect 20960 -3228 21056 -3212
rect 22372 -3212 22388 -2388
rect 22452 -3212 22468 -2388
rect 23784 -2388 23880 -2372
rect 22791 -2440 23513 -2439
rect 22791 -3160 22792 -2440
rect 23512 -3160 23513 -2440
rect 22791 -3161 23513 -3160
rect 22372 -3228 22468 -3212
rect 23784 -3212 23800 -2388
rect 23864 -3212 23880 -2388
rect 23784 -3228 23880 -3212
rect -22812 -3508 -22716 -3492
rect -23805 -3560 -23083 -3559
rect -23805 -4280 -23804 -3560
rect -23084 -4280 -23083 -3560
rect -23805 -4281 -23083 -4280
rect -22812 -4332 -22796 -3508
rect -22732 -4332 -22716 -3508
rect -21400 -3508 -21304 -3492
rect -22393 -3560 -21671 -3559
rect -22393 -4280 -22392 -3560
rect -21672 -4280 -21671 -3560
rect -22393 -4281 -21671 -4280
rect -22812 -4348 -22716 -4332
rect -21400 -4332 -21384 -3508
rect -21320 -4332 -21304 -3508
rect -19988 -3508 -19892 -3492
rect -20981 -3560 -20259 -3559
rect -20981 -4280 -20980 -3560
rect -20260 -4280 -20259 -3560
rect -20981 -4281 -20259 -4280
rect -21400 -4348 -21304 -4332
rect -19988 -4332 -19972 -3508
rect -19908 -4332 -19892 -3508
rect -18576 -3508 -18480 -3492
rect -19569 -3560 -18847 -3559
rect -19569 -4280 -19568 -3560
rect -18848 -4280 -18847 -3560
rect -19569 -4281 -18847 -4280
rect -19988 -4348 -19892 -4332
rect -18576 -4332 -18560 -3508
rect -18496 -4332 -18480 -3508
rect -17164 -3508 -17068 -3492
rect -18157 -3560 -17435 -3559
rect -18157 -4280 -18156 -3560
rect -17436 -4280 -17435 -3560
rect -18157 -4281 -17435 -4280
rect -18576 -4348 -18480 -4332
rect -17164 -4332 -17148 -3508
rect -17084 -4332 -17068 -3508
rect -15752 -3508 -15656 -3492
rect -16745 -3560 -16023 -3559
rect -16745 -4280 -16744 -3560
rect -16024 -4280 -16023 -3560
rect -16745 -4281 -16023 -4280
rect -17164 -4348 -17068 -4332
rect -15752 -4332 -15736 -3508
rect -15672 -4332 -15656 -3508
rect -14340 -3508 -14244 -3492
rect -15333 -3560 -14611 -3559
rect -15333 -4280 -15332 -3560
rect -14612 -4280 -14611 -3560
rect -15333 -4281 -14611 -4280
rect -15752 -4348 -15656 -4332
rect -14340 -4332 -14324 -3508
rect -14260 -4332 -14244 -3508
rect -12928 -3508 -12832 -3492
rect -13921 -3560 -13199 -3559
rect -13921 -4280 -13920 -3560
rect -13200 -4280 -13199 -3560
rect -13921 -4281 -13199 -4280
rect -14340 -4348 -14244 -4332
rect -12928 -4332 -12912 -3508
rect -12848 -4332 -12832 -3508
rect -11516 -3508 -11420 -3492
rect -12509 -3560 -11787 -3559
rect -12509 -4280 -12508 -3560
rect -11788 -4280 -11787 -3560
rect -12509 -4281 -11787 -4280
rect -12928 -4348 -12832 -4332
rect -11516 -4332 -11500 -3508
rect -11436 -4332 -11420 -3508
rect -10104 -3508 -10008 -3492
rect -11097 -3560 -10375 -3559
rect -11097 -4280 -11096 -3560
rect -10376 -4280 -10375 -3560
rect -11097 -4281 -10375 -4280
rect -11516 -4348 -11420 -4332
rect -10104 -4332 -10088 -3508
rect -10024 -4332 -10008 -3508
rect -8692 -3508 -8596 -3492
rect -9685 -3560 -8963 -3559
rect -9685 -4280 -9684 -3560
rect -8964 -4280 -8963 -3560
rect -9685 -4281 -8963 -4280
rect -10104 -4348 -10008 -4332
rect -8692 -4332 -8676 -3508
rect -8612 -4332 -8596 -3508
rect -7280 -3508 -7184 -3492
rect -8273 -3560 -7551 -3559
rect -8273 -4280 -8272 -3560
rect -7552 -4280 -7551 -3560
rect -8273 -4281 -7551 -4280
rect -8692 -4348 -8596 -4332
rect -7280 -4332 -7264 -3508
rect -7200 -4332 -7184 -3508
rect -5868 -3508 -5772 -3492
rect -6861 -3560 -6139 -3559
rect -6861 -4280 -6860 -3560
rect -6140 -4280 -6139 -3560
rect -6861 -4281 -6139 -4280
rect -7280 -4348 -7184 -4332
rect -5868 -4332 -5852 -3508
rect -5788 -4332 -5772 -3508
rect -4456 -3508 -4360 -3492
rect -5449 -3560 -4727 -3559
rect -5449 -4280 -5448 -3560
rect -4728 -4280 -4727 -3560
rect -5449 -4281 -4727 -4280
rect -5868 -4348 -5772 -4332
rect -4456 -4332 -4440 -3508
rect -4376 -4332 -4360 -3508
rect -3044 -3508 -2948 -3492
rect -4037 -3560 -3315 -3559
rect -4037 -4280 -4036 -3560
rect -3316 -4280 -3315 -3560
rect -4037 -4281 -3315 -4280
rect -4456 -4348 -4360 -4332
rect -3044 -4332 -3028 -3508
rect -2964 -4332 -2948 -3508
rect -1632 -3508 -1536 -3492
rect -2625 -3560 -1903 -3559
rect -2625 -4280 -2624 -3560
rect -1904 -4280 -1903 -3560
rect -2625 -4281 -1903 -4280
rect -3044 -4348 -2948 -4332
rect -1632 -4332 -1616 -3508
rect -1552 -4332 -1536 -3508
rect -220 -3508 -124 -3492
rect -1213 -3560 -491 -3559
rect -1213 -4280 -1212 -3560
rect -492 -4280 -491 -3560
rect -1213 -4281 -491 -4280
rect -1632 -4348 -1536 -4332
rect -220 -4332 -204 -3508
rect -140 -4332 -124 -3508
rect 1192 -3508 1288 -3492
rect 199 -3560 921 -3559
rect 199 -4280 200 -3560
rect 920 -4280 921 -3560
rect 199 -4281 921 -4280
rect -220 -4348 -124 -4332
rect 1192 -4332 1208 -3508
rect 1272 -4332 1288 -3508
rect 2604 -3508 2700 -3492
rect 1611 -3560 2333 -3559
rect 1611 -4280 1612 -3560
rect 2332 -4280 2333 -3560
rect 1611 -4281 2333 -4280
rect 1192 -4348 1288 -4332
rect 2604 -4332 2620 -3508
rect 2684 -4332 2700 -3508
rect 4016 -3508 4112 -3492
rect 3023 -3560 3745 -3559
rect 3023 -4280 3024 -3560
rect 3744 -4280 3745 -3560
rect 3023 -4281 3745 -4280
rect 2604 -4348 2700 -4332
rect 4016 -4332 4032 -3508
rect 4096 -4332 4112 -3508
rect 5428 -3508 5524 -3492
rect 4435 -3560 5157 -3559
rect 4435 -4280 4436 -3560
rect 5156 -4280 5157 -3560
rect 4435 -4281 5157 -4280
rect 4016 -4348 4112 -4332
rect 5428 -4332 5444 -3508
rect 5508 -4332 5524 -3508
rect 6840 -3508 6936 -3492
rect 5847 -3560 6569 -3559
rect 5847 -4280 5848 -3560
rect 6568 -4280 6569 -3560
rect 5847 -4281 6569 -4280
rect 5428 -4348 5524 -4332
rect 6840 -4332 6856 -3508
rect 6920 -4332 6936 -3508
rect 8252 -3508 8348 -3492
rect 7259 -3560 7981 -3559
rect 7259 -4280 7260 -3560
rect 7980 -4280 7981 -3560
rect 7259 -4281 7981 -4280
rect 6840 -4348 6936 -4332
rect 8252 -4332 8268 -3508
rect 8332 -4332 8348 -3508
rect 9664 -3508 9760 -3492
rect 8671 -3560 9393 -3559
rect 8671 -4280 8672 -3560
rect 9392 -4280 9393 -3560
rect 8671 -4281 9393 -4280
rect 8252 -4348 8348 -4332
rect 9664 -4332 9680 -3508
rect 9744 -4332 9760 -3508
rect 11076 -3508 11172 -3492
rect 10083 -3560 10805 -3559
rect 10083 -4280 10084 -3560
rect 10804 -4280 10805 -3560
rect 10083 -4281 10805 -4280
rect 9664 -4348 9760 -4332
rect 11076 -4332 11092 -3508
rect 11156 -4332 11172 -3508
rect 12488 -3508 12584 -3492
rect 11495 -3560 12217 -3559
rect 11495 -4280 11496 -3560
rect 12216 -4280 12217 -3560
rect 11495 -4281 12217 -4280
rect 11076 -4348 11172 -4332
rect 12488 -4332 12504 -3508
rect 12568 -4332 12584 -3508
rect 13900 -3508 13996 -3492
rect 12907 -3560 13629 -3559
rect 12907 -4280 12908 -3560
rect 13628 -4280 13629 -3560
rect 12907 -4281 13629 -4280
rect 12488 -4348 12584 -4332
rect 13900 -4332 13916 -3508
rect 13980 -4332 13996 -3508
rect 15312 -3508 15408 -3492
rect 14319 -3560 15041 -3559
rect 14319 -4280 14320 -3560
rect 15040 -4280 15041 -3560
rect 14319 -4281 15041 -4280
rect 13900 -4348 13996 -4332
rect 15312 -4332 15328 -3508
rect 15392 -4332 15408 -3508
rect 16724 -3508 16820 -3492
rect 15731 -3560 16453 -3559
rect 15731 -4280 15732 -3560
rect 16452 -4280 16453 -3560
rect 15731 -4281 16453 -4280
rect 15312 -4348 15408 -4332
rect 16724 -4332 16740 -3508
rect 16804 -4332 16820 -3508
rect 18136 -3508 18232 -3492
rect 17143 -3560 17865 -3559
rect 17143 -4280 17144 -3560
rect 17864 -4280 17865 -3560
rect 17143 -4281 17865 -4280
rect 16724 -4348 16820 -4332
rect 18136 -4332 18152 -3508
rect 18216 -4332 18232 -3508
rect 19548 -3508 19644 -3492
rect 18555 -3560 19277 -3559
rect 18555 -4280 18556 -3560
rect 19276 -4280 19277 -3560
rect 18555 -4281 19277 -4280
rect 18136 -4348 18232 -4332
rect 19548 -4332 19564 -3508
rect 19628 -4332 19644 -3508
rect 20960 -3508 21056 -3492
rect 19967 -3560 20689 -3559
rect 19967 -4280 19968 -3560
rect 20688 -4280 20689 -3560
rect 19967 -4281 20689 -4280
rect 19548 -4348 19644 -4332
rect 20960 -4332 20976 -3508
rect 21040 -4332 21056 -3508
rect 22372 -3508 22468 -3492
rect 21379 -3560 22101 -3559
rect 21379 -4280 21380 -3560
rect 22100 -4280 22101 -3560
rect 21379 -4281 22101 -4280
rect 20960 -4348 21056 -4332
rect 22372 -4332 22388 -3508
rect 22452 -4332 22468 -3508
rect 23784 -3508 23880 -3492
rect 22791 -3560 23513 -3559
rect 22791 -4280 22792 -3560
rect 23512 -4280 23513 -3560
rect 22791 -4281 23513 -4280
rect 22372 -4348 22468 -4332
rect 23784 -4332 23800 -3508
rect 23864 -4332 23880 -3508
rect 23784 -4348 23880 -4332
rect -22812 -4628 -22716 -4612
rect -23805 -4680 -23083 -4679
rect -23805 -5400 -23804 -4680
rect -23084 -5400 -23083 -4680
rect -23805 -5401 -23083 -5400
rect -22812 -5452 -22796 -4628
rect -22732 -5452 -22716 -4628
rect -21400 -4628 -21304 -4612
rect -22393 -4680 -21671 -4679
rect -22393 -5400 -22392 -4680
rect -21672 -5400 -21671 -4680
rect -22393 -5401 -21671 -5400
rect -22812 -5468 -22716 -5452
rect -21400 -5452 -21384 -4628
rect -21320 -5452 -21304 -4628
rect -19988 -4628 -19892 -4612
rect -20981 -4680 -20259 -4679
rect -20981 -5400 -20980 -4680
rect -20260 -5400 -20259 -4680
rect -20981 -5401 -20259 -5400
rect -21400 -5468 -21304 -5452
rect -19988 -5452 -19972 -4628
rect -19908 -5452 -19892 -4628
rect -18576 -4628 -18480 -4612
rect -19569 -4680 -18847 -4679
rect -19569 -5400 -19568 -4680
rect -18848 -5400 -18847 -4680
rect -19569 -5401 -18847 -5400
rect -19988 -5468 -19892 -5452
rect -18576 -5452 -18560 -4628
rect -18496 -5452 -18480 -4628
rect -17164 -4628 -17068 -4612
rect -18157 -4680 -17435 -4679
rect -18157 -5400 -18156 -4680
rect -17436 -5400 -17435 -4680
rect -18157 -5401 -17435 -5400
rect -18576 -5468 -18480 -5452
rect -17164 -5452 -17148 -4628
rect -17084 -5452 -17068 -4628
rect -15752 -4628 -15656 -4612
rect -16745 -4680 -16023 -4679
rect -16745 -5400 -16744 -4680
rect -16024 -5400 -16023 -4680
rect -16745 -5401 -16023 -5400
rect -17164 -5468 -17068 -5452
rect -15752 -5452 -15736 -4628
rect -15672 -5452 -15656 -4628
rect -14340 -4628 -14244 -4612
rect -15333 -4680 -14611 -4679
rect -15333 -5400 -15332 -4680
rect -14612 -5400 -14611 -4680
rect -15333 -5401 -14611 -5400
rect -15752 -5468 -15656 -5452
rect -14340 -5452 -14324 -4628
rect -14260 -5452 -14244 -4628
rect -12928 -4628 -12832 -4612
rect -13921 -4680 -13199 -4679
rect -13921 -5400 -13920 -4680
rect -13200 -5400 -13199 -4680
rect -13921 -5401 -13199 -5400
rect -14340 -5468 -14244 -5452
rect -12928 -5452 -12912 -4628
rect -12848 -5452 -12832 -4628
rect -11516 -4628 -11420 -4612
rect -12509 -4680 -11787 -4679
rect -12509 -5400 -12508 -4680
rect -11788 -5400 -11787 -4680
rect -12509 -5401 -11787 -5400
rect -12928 -5468 -12832 -5452
rect -11516 -5452 -11500 -4628
rect -11436 -5452 -11420 -4628
rect -10104 -4628 -10008 -4612
rect -11097 -4680 -10375 -4679
rect -11097 -5400 -11096 -4680
rect -10376 -5400 -10375 -4680
rect -11097 -5401 -10375 -5400
rect -11516 -5468 -11420 -5452
rect -10104 -5452 -10088 -4628
rect -10024 -5452 -10008 -4628
rect -8692 -4628 -8596 -4612
rect -9685 -4680 -8963 -4679
rect -9685 -5400 -9684 -4680
rect -8964 -5400 -8963 -4680
rect -9685 -5401 -8963 -5400
rect -10104 -5468 -10008 -5452
rect -8692 -5452 -8676 -4628
rect -8612 -5452 -8596 -4628
rect -7280 -4628 -7184 -4612
rect -8273 -4680 -7551 -4679
rect -8273 -5400 -8272 -4680
rect -7552 -5400 -7551 -4680
rect -8273 -5401 -7551 -5400
rect -8692 -5468 -8596 -5452
rect -7280 -5452 -7264 -4628
rect -7200 -5452 -7184 -4628
rect -5868 -4628 -5772 -4612
rect -6861 -4680 -6139 -4679
rect -6861 -5400 -6860 -4680
rect -6140 -5400 -6139 -4680
rect -6861 -5401 -6139 -5400
rect -7280 -5468 -7184 -5452
rect -5868 -5452 -5852 -4628
rect -5788 -5452 -5772 -4628
rect -4456 -4628 -4360 -4612
rect -5449 -4680 -4727 -4679
rect -5449 -5400 -5448 -4680
rect -4728 -5400 -4727 -4680
rect -5449 -5401 -4727 -5400
rect -5868 -5468 -5772 -5452
rect -4456 -5452 -4440 -4628
rect -4376 -5452 -4360 -4628
rect -3044 -4628 -2948 -4612
rect -4037 -4680 -3315 -4679
rect -4037 -5400 -4036 -4680
rect -3316 -5400 -3315 -4680
rect -4037 -5401 -3315 -5400
rect -4456 -5468 -4360 -5452
rect -3044 -5452 -3028 -4628
rect -2964 -5452 -2948 -4628
rect -1632 -4628 -1536 -4612
rect -2625 -4680 -1903 -4679
rect -2625 -5400 -2624 -4680
rect -1904 -5400 -1903 -4680
rect -2625 -5401 -1903 -5400
rect -3044 -5468 -2948 -5452
rect -1632 -5452 -1616 -4628
rect -1552 -5452 -1536 -4628
rect -220 -4628 -124 -4612
rect -1213 -4680 -491 -4679
rect -1213 -5400 -1212 -4680
rect -492 -5400 -491 -4680
rect -1213 -5401 -491 -5400
rect -1632 -5468 -1536 -5452
rect -220 -5452 -204 -4628
rect -140 -5452 -124 -4628
rect 1192 -4628 1288 -4612
rect 199 -4680 921 -4679
rect 199 -5400 200 -4680
rect 920 -5400 921 -4680
rect 199 -5401 921 -5400
rect -220 -5468 -124 -5452
rect 1192 -5452 1208 -4628
rect 1272 -5452 1288 -4628
rect 2604 -4628 2700 -4612
rect 1611 -4680 2333 -4679
rect 1611 -5400 1612 -4680
rect 2332 -5400 2333 -4680
rect 1611 -5401 2333 -5400
rect 1192 -5468 1288 -5452
rect 2604 -5452 2620 -4628
rect 2684 -5452 2700 -4628
rect 4016 -4628 4112 -4612
rect 3023 -4680 3745 -4679
rect 3023 -5400 3024 -4680
rect 3744 -5400 3745 -4680
rect 3023 -5401 3745 -5400
rect 2604 -5468 2700 -5452
rect 4016 -5452 4032 -4628
rect 4096 -5452 4112 -4628
rect 5428 -4628 5524 -4612
rect 4435 -4680 5157 -4679
rect 4435 -5400 4436 -4680
rect 5156 -5400 5157 -4680
rect 4435 -5401 5157 -5400
rect 4016 -5468 4112 -5452
rect 5428 -5452 5444 -4628
rect 5508 -5452 5524 -4628
rect 6840 -4628 6936 -4612
rect 5847 -4680 6569 -4679
rect 5847 -5400 5848 -4680
rect 6568 -5400 6569 -4680
rect 5847 -5401 6569 -5400
rect 5428 -5468 5524 -5452
rect 6840 -5452 6856 -4628
rect 6920 -5452 6936 -4628
rect 8252 -4628 8348 -4612
rect 7259 -4680 7981 -4679
rect 7259 -5400 7260 -4680
rect 7980 -5400 7981 -4680
rect 7259 -5401 7981 -5400
rect 6840 -5468 6936 -5452
rect 8252 -5452 8268 -4628
rect 8332 -5452 8348 -4628
rect 9664 -4628 9760 -4612
rect 8671 -4680 9393 -4679
rect 8671 -5400 8672 -4680
rect 9392 -5400 9393 -4680
rect 8671 -5401 9393 -5400
rect 8252 -5468 8348 -5452
rect 9664 -5452 9680 -4628
rect 9744 -5452 9760 -4628
rect 11076 -4628 11172 -4612
rect 10083 -4680 10805 -4679
rect 10083 -5400 10084 -4680
rect 10804 -5400 10805 -4680
rect 10083 -5401 10805 -5400
rect 9664 -5468 9760 -5452
rect 11076 -5452 11092 -4628
rect 11156 -5452 11172 -4628
rect 12488 -4628 12584 -4612
rect 11495 -4680 12217 -4679
rect 11495 -5400 11496 -4680
rect 12216 -5400 12217 -4680
rect 11495 -5401 12217 -5400
rect 11076 -5468 11172 -5452
rect 12488 -5452 12504 -4628
rect 12568 -5452 12584 -4628
rect 13900 -4628 13996 -4612
rect 12907 -4680 13629 -4679
rect 12907 -5400 12908 -4680
rect 13628 -5400 13629 -4680
rect 12907 -5401 13629 -5400
rect 12488 -5468 12584 -5452
rect 13900 -5452 13916 -4628
rect 13980 -5452 13996 -4628
rect 15312 -4628 15408 -4612
rect 14319 -4680 15041 -4679
rect 14319 -5400 14320 -4680
rect 15040 -5400 15041 -4680
rect 14319 -5401 15041 -5400
rect 13900 -5468 13996 -5452
rect 15312 -5452 15328 -4628
rect 15392 -5452 15408 -4628
rect 16724 -4628 16820 -4612
rect 15731 -4680 16453 -4679
rect 15731 -5400 15732 -4680
rect 16452 -5400 16453 -4680
rect 15731 -5401 16453 -5400
rect 15312 -5468 15408 -5452
rect 16724 -5452 16740 -4628
rect 16804 -5452 16820 -4628
rect 18136 -4628 18232 -4612
rect 17143 -4680 17865 -4679
rect 17143 -5400 17144 -4680
rect 17864 -5400 17865 -4680
rect 17143 -5401 17865 -5400
rect 16724 -5468 16820 -5452
rect 18136 -5452 18152 -4628
rect 18216 -5452 18232 -4628
rect 19548 -4628 19644 -4612
rect 18555 -4680 19277 -4679
rect 18555 -5400 18556 -4680
rect 19276 -5400 19277 -4680
rect 18555 -5401 19277 -5400
rect 18136 -5468 18232 -5452
rect 19548 -5452 19564 -4628
rect 19628 -5452 19644 -4628
rect 20960 -4628 21056 -4612
rect 19967 -4680 20689 -4679
rect 19967 -5400 19968 -4680
rect 20688 -5400 20689 -4680
rect 19967 -5401 20689 -5400
rect 19548 -5468 19644 -5452
rect 20960 -5452 20976 -4628
rect 21040 -5452 21056 -4628
rect 22372 -4628 22468 -4612
rect 21379 -4680 22101 -4679
rect 21379 -5400 21380 -4680
rect 22100 -5400 22101 -4680
rect 21379 -5401 22101 -5400
rect 20960 -5468 21056 -5452
rect 22372 -5452 22388 -4628
rect 22452 -5452 22468 -4628
rect 23784 -4628 23880 -4612
rect 22791 -4680 23513 -4679
rect 22791 -5400 22792 -4680
rect 23512 -5400 23513 -4680
rect 22791 -5401 23513 -5400
rect 22372 -5468 22468 -5452
rect 23784 -5452 23800 -4628
rect 23864 -5452 23880 -4628
rect 23784 -5468 23880 -5452
rect -22812 -5748 -22716 -5732
rect -23805 -5800 -23083 -5799
rect -23805 -6520 -23804 -5800
rect -23084 -6520 -23083 -5800
rect -23805 -6521 -23083 -6520
rect -22812 -6572 -22796 -5748
rect -22732 -6572 -22716 -5748
rect -21400 -5748 -21304 -5732
rect -22393 -5800 -21671 -5799
rect -22393 -6520 -22392 -5800
rect -21672 -6520 -21671 -5800
rect -22393 -6521 -21671 -6520
rect -22812 -6588 -22716 -6572
rect -21400 -6572 -21384 -5748
rect -21320 -6572 -21304 -5748
rect -19988 -5748 -19892 -5732
rect -20981 -5800 -20259 -5799
rect -20981 -6520 -20980 -5800
rect -20260 -6520 -20259 -5800
rect -20981 -6521 -20259 -6520
rect -21400 -6588 -21304 -6572
rect -19988 -6572 -19972 -5748
rect -19908 -6572 -19892 -5748
rect -18576 -5748 -18480 -5732
rect -19569 -5800 -18847 -5799
rect -19569 -6520 -19568 -5800
rect -18848 -6520 -18847 -5800
rect -19569 -6521 -18847 -6520
rect -19988 -6588 -19892 -6572
rect -18576 -6572 -18560 -5748
rect -18496 -6572 -18480 -5748
rect -17164 -5748 -17068 -5732
rect -18157 -5800 -17435 -5799
rect -18157 -6520 -18156 -5800
rect -17436 -6520 -17435 -5800
rect -18157 -6521 -17435 -6520
rect -18576 -6588 -18480 -6572
rect -17164 -6572 -17148 -5748
rect -17084 -6572 -17068 -5748
rect -15752 -5748 -15656 -5732
rect -16745 -5800 -16023 -5799
rect -16745 -6520 -16744 -5800
rect -16024 -6520 -16023 -5800
rect -16745 -6521 -16023 -6520
rect -17164 -6588 -17068 -6572
rect -15752 -6572 -15736 -5748
rect -15672 -6572 -15656 -5748
rect -14340 -5748 -14244 -5732
rect -15333 -5800 -14611 -5799
rect -15333 -6520 -15332 -5800
rect -14612 -6520 -14611 -5800
rect -15333 -6521 -14611 -6520
rect -15752 -6588 -15656 -6572
rect -14340 -6572 -14324 -5748
rect -14260 -6572 -14244 -5748
rect -12928 -5748 -12832 -5732
rect -13921 -5800 -13199 -5799
rect -13921 -6520 -13920 -5800
rect -13200 -6520 -13199 -5800
rect -13921 -6521 -13199 -6520
rect -14340 -6588 -14244 -6572
rect -12928 -6572 -12912 -5748
rect -12848 -6572 -12832 -5748
rect -11516 -5748 -11420 -5732
rect -12509 -5800 -11787 -5799
rect -12509 -6520 -12508 -5800
rect -11788 -6520 -11787 -5800
rect -12509 -6521 -11787 -6520
rect -12928 -6588 -12832 -6572
rect -11516 -6572 -11500 -5748
rect -11436 -6572 -11420 -5748
rect -10104 -5748 -10008 -5732
rect -11097 -5800 -10375 -5799
rect -11097 -6520 -11096 -5800
rect -10376 -6520 -10375 -5800
rect -11097 -6521 -10375 -6520
rect -11516 -6588 -11420 -6572
rect -10104 -6572 -10088 -5748
rect -10024 -6572 -10008 -5748
rect -8692 -5748 -8596 -5732
rect -9685 -5800 -8963 -5799
rect -9685 -6520 -9684 -5800
rect -8964 -6520 -8963 -5800
rect -9685 -6521 -8963 -6520
rect -10104 -6588 -10008 -6572
rect -8692 -6572 -8676 -5748
rect -8612 -6572 -8596 -5748
rect -7280 -5748 -7184 -5732
rect -8273 -5800 -7551 -5799
rect -8273 -6520 -8272 -5800
rect -7552 -6520 -7551 -5800
rect -8273 -6521 -7551 -6520
rect -8692 -6588 -8596 -6572
rect -7280 -6572 -7264 -5748
rect -7200 -6572 -7184 -5748
rect -5868 -5748 -5772 -5732
rect -6861 -5800 -6139 -5799
rect -6861 -6520 -6860 -5800
rect -6140 -6520 -6139 -5800
rect -6861 -6521 -6139 -6520
rect -7280 -6588 -7184 -6572
rect -5868 -6572 -5852 -5748
rect -5788 -6572 -5772 -5748
rect -4456 -5748 -4360 -5732
rect -5449 -5800 -4727 -5799
rect -5449 -6520 -5448 -5800
rect -4728 -6520 -4727 -5800
rect -5449 -6521 -4727 -6520
rect -5868 -6588 -5772 -6572
rect -4456 -6572 -4440 -5748
rect -4376 -6572 -4360 -5748
rect -3044 -5748 -2948 -5732
rect -4037 -5800 -3315 -5799
rect -4037 -6520 -4036 -5800
rect -3316 -6520 -3315 -5800
rect -4037 -6521 -3315 -6520
rect -4456 -6588 -4360 -6572
rect -3044 -6572 -3028 -5748
rect -2964 -6572 -2948 -5748
rect -1632 -5748 -1536 -5732
rect -2625 -5800 -1903 -5799
rect -2625 -6520 -2624 -5800
rect -1904 -6520 -1903 -5800
rect -2625 -6521 -1903 -6520
rect -3044 -6588 -2948 -6572
rect -1632 -6572 -1616 -5748
rect -1552 -6572 -1536 -5748
rect -220 -5748 -124 -5732
rect -1213 -5800 -491 -5799
rect -1213 -6520 -1212 -5800
rect -492 -6520 -491 -5800
rect -1213 -6521 -491 -6520
rect -1632 -6588 -1536 -6572
rect -220 -6572 -204 -5748
rect -140 -6572 -124 -5748
rect 1192 -5748 1288 -5732
rect 199 -5800 921 -5799
rect 199 -6520 200 -5800
rect 920 -6520 921 -5800
rect 199 -6521 921 -6520
rect -220 -6588 -124 -6572
rect 1192 -6572 1208 -5748
rect 1272 -6572 1288 -5748
rect 2604 -5748 2700 -5732
rect 1611 -5800 2333 -5799
rect 1611 -6520 1612 -5800
rect 2332 -6520 2333 -5800
rect 1611 -6521 2333 -6520
rect 1192 -6588 1288 -6572
rect 2604 -6572 2620 -5748
rect 2684 -6572 2700 -5748
rect 4016 -5748 4112 -5732
rect 3023 -5800 3745 -5799
rect 3023 -6520 3024 -5800
rect 3744 -6520 3745 -5800
rect 3023 -6521 3745 -6520
rect 2604 -6588 2700 -6572
rect 4016 -6572 4032 -5748
rect 4096 -6572 4112 -5748
rect 5428 -5748 5524 -5732
rect 4435 -5800 5157 -5799
rect 4435 -6520 4436 -5800
rect 5156 -6520 5157 -5800
rect 4435 -6521 5157 -6520
rect 4016 -6588 4112 -6572
rect 5428 -6572 5444 -5748
rect 5508 -6572 5524 -5748
rect 6840 -5748 6936 -5732
rect 5847 -5800 6569 -5799
rect 5847 -6520 5848 -5800
rect 6568 -6520 6569 -5800
rect 5847 -6521 6569 -6520
rect 5428 -6588 5524 -6572
rect 6840 -6572 6856 -5748
rect 6920 -6572 6936 -5748
rect 8252 -5748 8348 -5732
rect 7259 -5800 7981 -5799
rect 7259 -6520 7260 -5800
rect 7980 -6520 7981 -5800
rect 7259 -6521 7981 -6520
rect 6840 -6588 6936 -6572
rect 8252 -6572 8268 -5748
rect 8332 -6572 8348 -5748
rect 9664 -5748 9760 -5732
rect 8671 -5800 9393 -5799
rect 8671 -6520 8672 -5800
rect 9392 -6520 9393 -5800
rect 8671 -6521 9393 -6520
rect 8252 -6588 8348 -6572
rect 9664 -6572 9680 -5748
rect 9744 -6572 9760 -5748
rect 11076 -5748 11172 -5732
rect 10083 -5800 10805 -5799
rect 10083 -6520 10084 -5800
rect 10804 -6520 10805 -5800
rect 10083 -6521 10805 -6520
rect 9664 -6588 9760 -6572
rect 11076 -6572 11092 -5748
rect 11156 -6572 11172 -5748
rect 12488 -5748 12584 -5732
rect 11495 -5800 12217 -5799
rect 11495 -6520 11496 -5800
rect 12216 -6520 12217 -5800
rect 11495 -6521 12217 -6520
rect 11076 -6588 11172 -6572
rect 12488 -6572 12504 -5748
rect 12568 -6572 12584 -5748
rect 13900 -5748 13996 -5732
rect 12907 -5800 13629 -5799
rect 12907 -6520 12908 -5800
rect 13628 -6520 13629 -5800
rect 12907 -6521 13629 -6520
rect 12488 -6588 12584 -6572
rect 13900 -6572 13916 -5748
rect 13980 -6572 13996 -5748
rect 15312 -5748 15408 -5732
rect 14319 -5800 15041 -5799
rect 14319 -6520 14320 -5800
rect 15040 -6520 15041 -5800
rect 14319 -6521 15041 -6520
rect 13900 -6588 13996 -6572
rect 15312 -6572 15328 -5748
rect 15392 -6572 15408 -5748
rect 16724 -5748 16820 -5732
rect 15731 -5800 16453 -5799
rect 15731 -6520 15732 -5800
rect 16452 -6520 16453 -5800
rect 15731 -6521 16453 -6520
rect 15312 -6588 15408 -6572
rect 16724 -6572 16740 -5748
rect 16804 -6572 16820 -5748
rect 18136 -5748 18232 -5732
rect 17143 -5800 17865 -5799
rect 17143 -6520 17144 -5800
rect 17864 -6520 17865 -5800
rect 17143 -6521 17865 -6520
rect 16724 -6588 16820 -6572
rect 18136 -6572 18152 -5748
rect 18216 -6572 18232 -5748
rect 19548 -5748 19644 -5732
rect 18555 -5800 19277 -5799
rect 18555 -6520 18556 -5800
rect 19276 -6520 19277 -5800
rect 18555 -6521 19277 -6520
rect 18136 -6588 18232 -6572
rect 19548 -6572 19564 -5748
rect 19628 -6572 19644 -5748
rect 20960 -5748 21056 -5732
rect 19967 -5800 20689 -5799
rect 19967 -6520 19968 -5800
rect 20688 -6520 20689 -5800
rect 19967 -6521 20689 -6520
rect 19548 -6588 19644 -6572
rect 20960 -6572 20976 -5748
rect 21040 -6572 21056 -5748
rect 22372 -5748 22468 -5732
rect 21379 -5800 22101 -5799
rect 21379 -6520 21380 -5800
rect 22100 -6520 22101 -5800
rect 21379 -6521 22101 -6520
rect 20960 -6588 21056 -6572
rect 22372 -6572 22388 -5748
rect 22452 -6572 22468 -5748
rect 23784 -5748 23880 -5732
rect 22791 -5800 23513 -5799
rect 22791 -6520 22792 -5800
rect 23512 -6520 23513 -5800
rect 22791 -6521 23513 -6520
rect 22372 -6588 22468 -6572
rect 23784 -6572 23800 -5748
rect 23864 -6572 23880 -5748
rect 23784 -6588 23880 -6572
rect -22812 -6868 -22716 -6852
rect -23805 -6920 -23083 -6919
rect -23805 -7640 -23804 -6920
rect -23084 -7640 -23083 -6920
rect -23805 -7641 -23083 -7640
rect -22812 -7692 -22796 -6868
rect -22732 -7692 -22716 -6868
rect -21400 -6868 -21304 -6852
rect -22393 -6920 -21671 -6919
rect -22393 -7640 -22392 -6920
rect -21672 -7640 -21671 -6920
rect -22393 -7641 -21671 -7640
rect -22812 -7708 -22716 -7692
rect -21400 -7692 -21384 -6868
rect -21320 -7692 -21304 -6868
rect -19988 -6868 -19892 -6852
rect -20981 -6920 -20259 -6919
rect -20981 -7640 -20980 -6920
rect -20260 -7640 -20259 -6920
rect -20981 -7641 -20259 -7640
rect -21400 -7708 -21304 -7692
rect -19988 -7692 -19972 -6868
rect -19908 -7692 -19892 -6868
rect -18576 -6868 -18480 -6852
rect -19569 -6920 -18847 -6919
rect -19569 -7640 -19568 -6920
rect -18848 -7640 -18847 -6920
rect -19569 -7641 -18847 -7640
rect -19988 -7708 -19892 -7692
rect -18576 -7692 -18560 -6868
rect -18496 -7692 -18480 -6868
rect -17164 -6868 -17068 -6852
rect -18157 -6920 -17435 -6919
rect -18157 -7640 -18156 -6920
rect -17436 -7640 -17435 -6920
rect -18157 -7641 -17435 -7640
rect -18576 -7708 -18480 -7692
rect -17164 -7692 -17148 -6868
rect -17084 -7692 -17068 -6868
rect -15752 -6868 -15656 -6852
rect -16745 -6920 -16023 -6919
rect -16745 -7640 -16744 -6920
rect -16024 -7640 -16023 -6920
rect -16745 -7641 -16023 -7640
rect -17164 -7708 -17068 -7692
rect -15752 -7692 -15736 -6868
rect -15672 -7692 -15656 -6868
rect -14340 -6868 -14244 -6852
rect -15333 -6920 -14611 -6919
rect -15333 -7640 -15332 -6920
rect -14612 -7640 -14611 -6920
rect -15333 -7641 -14611 -7640
rect -15752 -7708 -15656 -7692
rect -14340 -7692 -14324 -6868
rect -14260 -7692 -14244 -6868
rect -12928 -6868 -12832 -6852
rect -13921 -6920 -13199 -6919
rect -13921 -7640 -13920 -6920
rect -13200 -7640 -13199 -6920
rect -13921 -7641 -13199 -7640
rect -14340 -7708 -14244 -7692
rect -12928 -7692 -12912 -6868
rect -12848 -7692 -12832 -6868
rect -11516 -6868 -11420 -6852
rect -12509 -6920 -11787 -6919
rect -12509 -7640 -12508 -6920
rect -11788 -7640 -11787 -6920
rect -12509 -7641 -11787 -7640
rect -12928 -7708 -12832 -7692
rect -11516 -7692 -11500 -6868
rect -11436 -7692 -11420 -6868
rect -10104 -6868 -10008 -6852
rect -11097 -6920 -10375 -6919
rect -11097 -7640 -11096 -6920
rect -10376 -7640 -10375 -6920
rect -11097 -7641 -10375 -7640
rect -11516 -7708 -11420 -7692
rect -10104 -7692 -10088 -6868
rect -10024 -7692 -10008 -6868
rect -8692 -6868 -8596 -6852
rect -9685 -6920 -8963 -6919
rect -9685 -7640 -9684 -6920
rect -8964 -7640 -8963 -6920
rect -9685 -7641 -8963 -7640
rect -10104 -7708 -10008 -7692
rect -8692 -7692 -8676 -6868
rect -8612 -7692 -8596 -6868
rect -7280 -6868 -7184 -6852
rect -8273 -6920 -7551 -6919
rect -8273 -7640 -8272 -6920
rect -7552 -7640 -7551 -6920
rect -8273 -7641 -7551 -7640
rect -8692 -7708 -8596 -7692
rect -7280 -7692 -7264 -6868
rect -7200 -7692 -7184 -6868
rect -5868 -6868 -5772 -6852
rect -6861 -6920 -6139 -6919
rect -6861 -7640 -6860 -6920
rect -6140 -7640 -6139 -6920
rect -6861 -7641 -6139 -7640
rect -7280 -7708 -7184 -7692
rect -5868 -7692 -5852 -6868
rect -5788 -7692 -5772 -6868
rect -4456 -6868 -4360 -6852
rect -5449 -6920 -4727 -6919
rect -5449 -7640 -5448 -6920
rect -4728 -7640 -4727 -6920
rect -5449 -7641 -4727 -7640
rect -5868 -7708 -5772 -7692
rect -4456 -7692 -4440 -6868
rect -4376 -7692 -4360 -6868
rect -3044 -6868 -2948 -6852
rect -4037 -6920 -3315 -6919
rect -4037 -7640 -4036 -6920
rect -3316 -7640 -3315 -6920
rect -4037 -7641 -3315 -7640
rect -4456 -7708 -4360 -7692
rect -3044 -7692 -3028 -6868
rect -2964 -7692 -2948 -6868
rect -1632 -6868 -1536 -6852
rect -2625 -6920 -1903 -6919
rect -2625 -7640 -2624 -6920
rect -1904 -7640 -1903 -6920
rect -2625 -7641 -1903 -7640
rect -3044 -7708 -2948 -7692
rect -1632 -7692 -1616 -6868
rect -1552 -7692 -1536 -6868
rect -220 -6868 -124 -6852
rect -1213 -6920 -491 -6919
rect -1213 -7640 -1212 -6920
rect -492 -7640 -491 -6920
rect -1213 -7641 -491 -7640
rect -1632 -7708 -1536 -7692
rect -220 -7692 -204 -6868
rect -140 -7692 -124 -6868
rect 1192 -6868 1288 -6852
rect 199 -6920 921 -6919
rect 199 -7640 200 -6920
rect 920 -7640 921 -6920
rect 199 -7641 921 -7640
rect -220 -7708 -124 -7692
rect 1192 -7692 1208 -6868
rect 1272 -7692 1288 -6868
rect 2604 -6868 2700 -6852
rect 1611 -6920 2333 -6919
rect 1611 -7640 1612 -6920
rect 2332 -7640 2333 -6920
rect 1611 -7641 2333 -7640
rect 1192 -7708 1288 -7692
rect 2604 -7692 2620 -6868
rect 2684 -7692 2700 -6868
rect 4016 -6868 4112 -6852
rect 3023 -6920 3745 -6919
rect 3023 -7640 3024 -6920
rect 3744 -7640 3745 -6920
rect 3023 -7641 3745 -7640
rect 2604 -7708 2700 -7692
rect 4016 -7692 4032 -6868
rect 4096 -7692 4112 -6868
rect 5428 -6868 5524 -6852
rect 4435 -6920 5157 -6919
rect 4435 -7640 4436 -6920
rect 5156 -7640 5157 -6920
rect 4435 -7641 5157 -7640
rect 4016 -7708 4112 -7692
rect 5428 -7692 5444 -6868
rect 5508 -7692 5524 -6868
rect 6840 -6868 6936 -6852
rect 5847 -6920 6569 -6919
rect 5847 -7640 5848 -6920
rect 6568 -7640 6569 -6920
rect 5847 -7641 6569 -7640
rect 5428 -7708 5524 -7692
rect 6840 -7692 6856 -6868
rect 6920 -7692 6936 -6868
rect 8252 -6868 8348 -6852
rect 7259 -6920 7981 -6919
rect 7259 -7640 7260 -6920
rect 7980 -7640 7981 -6920
rect 7259 -7641 7981 -7640
rect 6840 -7708 6936 -7692
rect 8252 -7692 8268 -6868
rect 8332 -7692 8348 -6868
rect 9664 -6868 9760 -6852
rect 8671 -6920 9393 -6919
rect 8671 -7640 8672 -6920
rect 9392 -7640 9393 -6920
rect 8671 -7641 9393 -7640
rect 8252 -7708 8348 -7692
rect 9664 -7692 9680 -6868
rect 9744 -7692 9760 -6868
rect 11076 -6868 11172 -6852
rect 10083 -6920 10805 -6919
rect 10083 -7640 10084 -6920
rect 10804 -7640 10805 -6920
rect 10083 -7641 10805 -7640
rect 9664 -7708 9760 -7692
rect 11076 -7692 11092 -6868
rect 11156 -7692 11172 -6868
rect 12488 -6868 12584 -6852
rect 11495 -6920 12217 -6919
rect 11495 -7640 11496 -6920
rect 12216 -7640 12217 -6920
rect 11495 -7641 12217 -7640
rect 11076 -7708 11172 -7692
rect 12488 -7692 12504 -6868
rect 12568 -7692 12584 -6868
rect 13900 -6868 13996 -6852
rect 12907 -6920 13629 -6919
rect 12907 -7640 12908 -6920
rect 13628 -7640 13629 -6920
rect 12907 -7641 13629 -7640
rect 12488 -7708 12584 -7692
rect 13900 -7692 13916 -6868
rect 13980 -7692 13996 -6868
rect 15312 -6868 15408 -6852
rect 14319 -6920 15041 -6919
rect 14319 -7640 14320 -6920
rect 15040 -7640 15041 -6920
rect 14319 -7641 15041 -7640
rect 13900 -7708 13996 -7692
rect 15312 -7692 15328 -6868
rect 15392 -7692 15408 -6868
rect 16724 -6868 16820 -6852
rect 15731 -6920 16453 -6919
rect 15731 -7640 15732 -6920
rect 16452 -7640 16453 -6920
rect 15731 -7641 16453 -7640
rect 15312 -7708 15408 -7692
rect 16724 -7692 16740 -6868
rect 16804 -7692 16820 -6868
rect 18136 -6868 18232 -6852
rect 17143 -6920 17865 -6919
rect 17143 -7640 17144 -6920
rect 17864 -7640 17865 -6920
rect 17143 -7641 17865 -7640
rect 16724 -7708 16820 -7692
rect 18136 -7692 18152 -6868
rect 18216 -7692 18232 -6868
rect 19548 -6868 19644 -6852
rect 18555 -6920 19277 -6919
rect 18555 -7640 18556 -6920
rect 19276 -7640 19277 -6920
rect 18555 -7641 19277 -7640
rect 18136 -7708 18232 -7692
rect 19548 -7692 19564 -6868
rect 19628 -7692 19644 -6868
rect 20960 -6868 21056 -6852
rect 19967 -6920 20689 -6919
rect 19967 -7640 19968 -6920
rect 20688 -7640 20689 -6920
rect 19967 -7641 20689 -7640
rect 19548 -7708 19644 -7692
rect 20960 -7692 20976 -6868
rect 21040 -7692 21056 -6868
rect 22372 -6868 22468 -6852
rect 21379 -6920 22101 -6919
rect 21379 -7640 21380 -6920
rect 22100 -7640 22101 -6920
rect 21379 -7641 22101 -7640
rect 20960 -7708 21056 -7692
rect 22372 -7692 22388 -6868
rect 22452 -7692 22468 -6868
rect 23784 -6868 23880 -6852
rect 22791 -6920 23513 -6919
rect 22791 -7640 22792 -6920
rect 23512 -7640 23513 -6920
rect 22791 -7641 23513 -7640
rect 22372 -7708 22468 -7692
rect 23784 -7692 23800 -6868
rect 23864 -7692 23880 -6868
rect 23784 -7708 23880 -7692
rect -22812 -7988 -22716 -7972
rect -23805 -8040 -23083 -8039
rect -23805 -8760 -23804 -8040
rect -23084 -8760 -23083 -8040
rect -23805 -8761 -23083 -8760
rect -22812 -8812 -22796 -7988
rect -22732 -8812 -22716 -7988
rect -21400 -7988 -21304 -7972
rect -22393 -8040 -21671 -8039
rect -22393 -8760 -22392 -8040
rect -21672 -8760 -21671 -8040
rect -22393 -8761 -21671 -8760
rect -22812 -8828 -22716 -8812
rect -21400 -8812 -21384 -7988
rect -21320 -8812 -21304 -7988
rect -19988 -7988 -19892 -7972
rect -20981 -8040 -20259 -8039
rect -20981 -8760 -20980 -8040
rect -20260 -8760 -20259 -8040
rect -20981 -8761 -20259 -8760
rect -21400 -8828 -21304 -8812
rect -19988 -8812 -19972 -7988
rect -19908 -8812 -19892 -7988
rect -18576 -7988 -18480 -7972
rect -19569 -8040 -18847 -8039
rect -19569 -8760 -19568 -8040
rect -18848 -8760 -18847 -8040
rect -19569 -8761 -18847 -8760
rect -19988 -8828 -19892 -8812
rect -18576 -8812 -18560 -7988
rect -18496 -8812 -18480 -7988
rect -17164 -7988 -17068 -7972
rect -18157 -8040 -17435 -8039
rect -18157 -8760 -18156 -8040
rect -17436 -8760 -17435 -8040
rect -18157 -8761 -17435 -8760
rect -18576 -8828 -18480 -8812
rect -17164 -8812 -17148 -7988
rect -17084 -8812 -17068 -7988
rect -15752 -7988 -15656 -7972
rect -16745 -8040 -16023 -8039
rect -16745 -8760 -16744 -8040
rect -16024 -8760 -16023 -8040
rect -16745 -8761 -16023 -8760
rect -17164 -8828 -17068 -8812
rect -15752 -8812 -15736 -7988
rect -15672 -8812 -15656 -7988
rect -14340 -7988 -14244 -7972
rect -15333 -8040 -14611 -8039
rect -15333 -8760 -15332 -8040
rect -14612 -8760 -14611 -8040
rect -15333 -8761 -14611 -8760
rect -15752 -8828 -15656 -8812
rect -14340 -8812 -14324 -7988
rect -14260 -8812 -14244 -7988
rect -12928 -7988 -12832 -7972
rect -13921 -8040 -13199 -8039
rect -13921 -8760 -13920 -8040
rect -13200 -8760 -13199 -8040
rect -13921 -8761 -13199 -8760
rect -14340 -8828 -14244 -8812
rect -12928 -8812 -12912 -7988
rect -12848 -8812 -12832 -7988
rect -11516 -7988 -11420 -7972
rect -12509 -8040 -11787 -8039
rect -12509 -8760 -12508 -8040
rect -11788 -8760 -11787 -8040
rect -12509 -8761 -11787 -8760
rect -12928 -8828 -12832 -8812
rect -11516 -8812 -11500 -7988
rect -11436 -8812 -11420 -7988
rect -10104 -7988 -10008 -7972
rect -11097 -8040 -10375 -8039
rect -11097 -8760 -11096 -8040
rect -10376 -8760 -10375 -8040
rect -11097 -8761 -10375 -8760
rect -11516 -8828 -11420 -8812
rect -10104 -8812 -10088 -7988
rect -10024 -8812 -10008 -7988
rect -8692 -7988 -8596 -7972
rect -9685 -8040 -8963 -8039
rect -9685 -8760 -9684 -8040
rect -8964 -8760 -8963 -8040
rect -9685 -8761 -8963 -8760
rect -10104 -8828 -10008 -8812
rect -8692 -8812 -8676 -7988
rect -8612 -8812 -8596 -7988
rect -7280 -7988 -7184 -7972
rect -8273 -8040 -7551 -8039
rect -8273 -8760 -8272 -8040
rect -7552 -8760 -7551 -8040
rect -8273 -8761 -7551 -8760
rect -8692 -8828 -8596 -8812
rect -7280 -8812 -7264 -7988
rect -7200 -8812 -7184 -7988
rect -5868 -7988 -5772 -7972
rect -6861 -8040 -6139 -8039
rect -6861 -8760 -6860 -8040
rect -6140 -8760 -6139 -8040
rect -6861 -8761 -6139 -8760
rect -7280 -8828 -7184 -8812
rect -5868 -8812 -5852 -7988
rect -5788 -8812 -5772 -7988
rect -4456 -7988 -4360 -7972
rect -5449 -8040 -4727 -8039
rect -5449 -8760 -5448 -8040
rect -4728 -8760 -4727 -8040
rect -5449 -8761 -4727 -8760
rect -5868 -8828 -5772 -8812
rect -4456 -8812 -4440 -7988
rect -4376 -8812 -4360 -7988
rect -3044 -7988 -2948 -7972
rect -4037 -8040 -3315 -8039
rect -4037 -8760 -4036 -8040
rect -3316 -8760 -3315 -8040
rect -4037 -8761 -3315 -8760
rect -4456 -8828 -4360 -8812
rect -3044 -8812 -3028 -7988
rect -2964 -8812 -2948 -7988
rect -1632 -7988 -1536 -7972
rect -2625 -8040 -1903 -8039
rect -2625 -8760 -2624 -8040
rect -1904 -8760 -1903 -8040
rect -2625 -8761 -1903 -8760
rect -3044 -8828 -2948 -8812
rect -1632 -8812 -1616 -7988
rect -1552 -8812 -1536 -7988
rect -220 -7988 -124 -7972
rect -1213 -8040 -491 -8039
rect -1213 -8760 -1212 -8040
rect -492 -8760 -491 -8040
rect -1213 -8761 -491 -8760
rect -1632 -8828 -1536 -8812
rect -220 -8812 -204 -7988
rect -140 -8812 -124 -7988
rect 1192 -7988 1288 -7972
rect 199 -8040 921 -8039
rect 199 -8760 200 -8040
rect 920 -8760 921 -8040
rect 199 -8761 921 -8760
rect -220 -8828 -124 -8812
rect 1192 -8812 1208 -7988
rect 1272 -8812 1288 -7988
rect 2604 -7988 2700 -7972
rect 1611 -8040 2333 -8039
rect 1611 -8760 1612 -8040
rect 2332 -8760 2333 -8040
rect 1611 -8761 2333 -8760
rect 1192 -8828 1288 -8812
rect 2604 -8812 2620 -7988
rect 2684 -8812 2700 -7988
rect 4016 -7988 4112 -7972
rect 3023 -8040 3745 -8039
rect 3023 -8760 3024 -8040
rect 3744 -8760 3745 -8040
rect 3023 -8761 3745 -8760
rect 2604 -8828 2700 -8812
rect 4016 -8812 4032 -7988
rect 4096 -8812 4112 -7988
rect 5428 -7988 5524 -7972
rect 4435 -8040 5157 -8039
rect 4435 -8760 4436 -8040
rect 5156 -8760 5157 -8040
rect 4435 -8761 5157 -8760
rect 4016 -8828 4112 -8812
rect 5428 -8812 5444 -7988
rect 5508 -8812 5524 -7988
rect 6840 -7988 6936 -7972
rect 5847 -8040 6569 -8039
rect 5847 -8760 5848 -8040
rect 6568 -8760 6569 -8040
rect 5847 -8761 6569 -8760
rect 5428 -8828 5524 -8812
rect 6840 -8812 6856 -7988
rect 6920 -8812 6936 -7988
rect 8252 -7988 8348 -7972
rect 7259 -8040 7981 -8039
rect 7259 -8760 7260 -8040
rect 7980 -8760 7981 -8040
rect 7259 -8761 7981 -8760
rect 6840 -8828 6936 -8812
rect 8252 -8812 8268 -7988
rect 8332 -8812 8348 -7988
rect 9664 -7988 9760 -7972
rect 8671 -8040 9393 -8039
rect 8671 -8760 8672 -8040
rect 9392 -8760 9393 -8040
rect 8671 -8761 9393 -8760
rect 8252 -8828 8348 -8812
rect 9664 -8812 9680 -7988
rect 9744 -8812 9760 -7988
rect 11076 -7988 11172 -7972
rect 10083 -8040 10805 -8039
rect 10083 -8760 10084 -8040
rect 10804 -8760 10805 -8040
rect 10083 -8761 10805 -8760
rect 9664 -8828 9760 -8812
rect 11076 -8812 11092 -7988
rect 11156 -8812 11172 -7988
rect 12488 -7988 12584 -7972
rect 11495 -8040 12217 -8039
rect 11495 -8760 11496 -8040
rect 12216 -8760 12217 -8040
rect 11495 -8761 12217 -8760
rect 11076 -8828 11172 -8812
rect 12488 -8812 12504 -7988
rect 12568 -8812 12584 -7988
rect 13900 -7988 13996 -7972
rect 12907 -8040 13629 -8039
rect 12907 -8760 12908 -8040
rect 13628 -8760 13629 -8040
rect 12907 -8761 13629 -8760
rect 12488 -8828 12584 -8812
rect 13900 -8812 13916 -7988
rect 13980 -8812 13996 -7988
rect 15312 -7988 15408 -7972
rect 14319 -8040 15041 -8039
rect 14319 -8760 14320 -8040
rect 15040 -8760 15041 -8040
rect 14319 -8761 15041 -8760
rect 13900 -8828 13996 -8812
rect 15312 -8812 15328 -7988
rect 15392 -8812 15408 -7988
rect 16724 -7988 16820 -7972
rect 15731 -8040 16453 -8039
rect 15731 -8760 15732 -8040
rect 16452 -8760 16453 -8040
rect 15731 -8761 16453 -8760
rect 15312 -8828 15408 -8812
rect 16724 -8812 16740 -7988
rect 16804 -8812 16820 -7988
rect 18136 -7988 18232 -7972
rect 17143 -8040 17865 -8039
rect 17143 -8760 17144 -8040
rect 17864 -8760 17865 -8040
rect 17143 -8761 17865 -8760
rect 16724 -8828 16820 -8812
rect 18136 -8812 18152 -7988
rect 18216 -8812 18232 -7988
rect 19548 -7988 19644 -7972
rect 18555 -8040 19277 -8039
rect 18555 -8760 18556 -8040
rect 19276 -8760 19277 -8040
rect 18555 -8761 19277 -8760
rect 18136 -8828 18232 -8812
rect 19548 -8812 19564 -7988
rect 19628 -8812 19644 -7988
rect 20960 -7988 21056 -7972
rect 19967 -8040 20689 -8039
rect 19967 -8760 19968 -8040
rect 20688 -8760 20689 -8040
rect 19967 -8761 20689 -8760
rect 19548 -8828 19644 -8812
rect 20960 -8812 20976 -7988
rect 21040 -8812 21056 -7988
rect 22372 -7988 22468 -7972
rect 21379 -8040 22101 -8039
rect 21379 -8760 21380 -8040
rect 22100 -8760 22101 -8040
rect 21379 -8761 22101 -8760
rect 20960 -8828 21056 -8812
rect 22372 -8812 22388 -7988
rect 22452 -8812 22468 -7988
rect 23784 -7988 23880 -7972
rect 22791 -8040 23513 -8039
rect 22791 -8760 22792 -8040
rect 23512 -8760 23513 -8040
rect 22791 -8761 23513 -8760
rect 22372 -8828 22468 -8812
rect 23784 -8812 23800 -7988
rect 23864 -8812 23880 -7988
rect 23784 -8828 23880 -8812
rect -22812 -9108 -22716 -9092
rect -23805 -9160 -23083 -9159
rect -23805 -9880 -23804 -9160
rect -23084 -9880 -23083 -9160
rect -23805 -9881 -23083 -9880
rect -22812 -9932 -22796 -9108
rect -22732 -9932 -22716 -9108
rect -21400 -9108 -21304 -9092
rect -22393 -9160 -21671 -9159
rect -22393 -9880 -22392 -9160
rect -21672 -9880 -21671 -9160
rect -22393 -9881 -21671 -9880
rect -22812 -9948 -22716 -9932
rect -21400 -9932 -21384 -9108
rect -21320 -9932 -21304 -9108
rect -19988 -9108 -19892 -9092
rect -20981 -9160 -20259 -9159
rect -20981 -9880 -20980 -9160
rect -20260 -9880 -20259 -9160
rect -20981 -9881 -20259 -9880
rect -21400 -9948 -21304 -9932
rect -19988 -9932 -19972 -9108
rect -19908 -9932 -19892 -9108
rect -18576 -9108 -18480 -9092
rect -19569 -9160 -18847 -9159
rect -19569 -9880 -19568 -9160
rect -18848 -9880 -18847 -9160
rect -19569 -9881 -18847 -9880
rect -19988 -9948 -19892 -9932
rect -18576 -9932 -18560 -9108
rect -18496 -9932 -18480 -9108
rect -17164 -9108 -17068 -9092
rect -18157 -9160 -17435 -9159
rect -18157 -9880 -18156 -9160
rect -17436 -9880 -17435 -9160
rect -18157 -9881 -17435 -9880
rect -18576 -9948 -18480 -9932
rect -17164 -9932 -17148 -9108
rect -17084 -9932 -17068 -9108
rect -15752 -9108 -15656 -9092
rect -16745 -9160 -16023 -9159
rect -16745 -9880 -16744 -9160
rect -16024 -9880 -16023 -9160
rect -16745 -9881 -16023 -9880
rect -17164 -9948 -17068 -9932
rect -15752 -9932 -15736 -9108
rect -15672 -9932 -15656 -9108
rect -14340 -9108 -14244 -9092
rect -15333 -9160 -14611 -9159
rect -15333 -9880 -15332 -9160
rect -14612 -9880 -14611 -9160
rect -15333 -9881 -14611 -9880
rect -15752 -9948 -15656 -9932
rect -14340 -9932 -14324 -9108
rect -14260 -9932 -14244 -9108
rect -12928 -9108 -12832 -9092
rect -13921 -9160 -13199 -9159
rect -13921 -9880 -13920 -9160
rect -13200 -9880 -13199 -9160
rect -13921 -9881 -13199 -9880
rect -14340 -9948 -14244 -9932
rect -12928 -9932 -12912 -9108
rect -12848 -9932 -12832 -9108
rect -11516 -9108 -11420 -9092
rect -12509 -9160 -11787 -9159
rect -12509 -9880 -12508 -9160
rect -11788 -9880 -11787 -9160
rect -12509 -9881 -11787 -9880
rect -12928 -9948 -12832 -9932
rect -11516 -9932 -11500 -9108
rect -11436 -9932 -11420 -9108
rect -10104 -9108 -10008 -9092
rect -11097 -9160 -10375 -9159
rect -11097 -9880 -11096 -9160
rect -10376 -9880 -10375 -9160
rect -11097 -9881 -10375 -9880
rect -11516 -9948 -11420 -9932
rect -10104 -9932 -10088 -9108
rect -10024 -9932 -10008 -9108
rect -8692 -9108 -8596 -9092
rect -9685 -9160 -8963 -9159
rect -9685 -9880 -9684 -9160
rect -8964 -9880 -8963 -9160
rect -9685 -9881 -8963 -9880
rect -10104 -9948 -10008 -9932
rect -8692 -9932 -8676 -9108
rect -8612 -9932 -8596 -9108
rect -7280 -9108 -7184 -9092
rect -8273 -9160 -7551 -9159
rect -8273 -9880 -8272 -9160
rect -7552 -9880 -7551 -9160
rect -8273 -9881 -7551 -9880
rect -8692 -9948 -8596 -9932
rect -7280 -9932 -7264 -9108
rect -7200 -9932 -7184 -9108
rect -5868 -9108 -5772 -9092
rect -6861 -9160 -6139 -9159
rect -6861 -9880 -6860 -9160
rect -6140 -9880 -6139 -9160
rect -6861 -9881 -6139 -9880
rect -7280 -9948 -7184 -9932
rect -5868 -9932 -5852 -9108
rect -5788 -9932 -5772 -9108
rect -4456 -9108 -4360 -9092
rect -5449 -9160 -4727 -9159
rect -5449 -9880 -5448 -9160
rect -4728 -9880 -4727 -9160
rect -5449 -9881 -4727 -9880
rect -5868 -9948 -5772 -9932
rect -4456 -9932 -4440 -9108
rect -4376 -9932 -4360 -9108
rect -3044 -9108 -2948 -9092
rect -4037 -9160 -3315 -9159
rect -4037 -9880 -4036 -9160
rect -3316 -9880 -3315 -9160
rect -4037 -9881 -3315 -9880
rect -4456 -9948 -4360 -9932
rect -3044 -9932 -3028 -9108
rect -2964 -9932 -2948 -9108
rect -1632 -9108 -1536 -9092
rect -2625 -9160 -1903 -9159
rect -2625 -9880 -2624 -9160
rect -1904 -9880 -1903 -9160
rect -2625 -9881 -1903 -9880
rect -3044 -9948 -2948 -9932
rect -1632 -9932 -1616 -9108
rect -1552 -9932 -1536 -9108
rect -220 -9108 -124 -9092
rect -1213 -9160 -491 -9159
rect -1213 -9880 -1212 -9160
rect -492 -9880 -491 -9160
rect -1213 -9881 -491 -9880
rect -1632 -9948 -1536 -9932
rect -220 -9932 -204 -9108
rect -140 -9932 -124 -9108
rect 1192 -9108 1288 -9092
rect 199 -9160 921 -9159
rect 199 -9880 200 -9160
rect 920 -9880 921 -9160
rect 199 -9881 921 -9880
rect -220 -9948 -124 -9932
rect 1192 -9932 1208 -9108
rect 1272 -9932 1288 -9108
rect 2604 -9108 2700 -9092
rect 1611 -9160 2333 -9159
rect 1611 -9880 1612 -9160
rect 2332 -9880 2333 -9160
rect 1611 -9881 2333 -9880
rect 1192 -9948 1288 -9932
rect 2604 -9932 2620 -9108
rect 2684 -9932 2700 -9108
rect 4016 -9108 4112 -9092
rect 3023 -9160 3745 -9159
rect 3023 -9880 3024 -9160
rect 3744 -9880 3745 -9160
rect 3023 -9881 3745 -9880
rect 2604 -9948 2700 -9932
rect 4016 -9932 4032 -9108
rect 4096 -9932 4112 -9108
rect 5428 -9108 5524 -9092
rect 4435 -9160 5157 -9159
rect 4435 -9880 4436 -9160
rect 5156 -9880 5157 -9160
rect 4435 -9881 5157 -9880
rect 4016 -9948 4112 -9932
rect 5428 -9932 5444 -9108
rect 5508 -9932 5524 -9108
rect 6840 -9108 6936 -9092
rect 5847 -9160 6569 -9159
rect 5847 -9880 5848 -9160
rect 6568 -9880 6569 -9160
rect 5847 -9881 6569 -9880
rect 5428 -9948 5524 -9932
rect 6840 -9932 6856 -9108
rect 6920 -9932 6936 -9108
rect 8252 -9108 8348 -9092
rect 7259 -9160 7981 -9159
rect 7259 -9880 7260 -9160
rect 7980 -9880 7981 -9160
rect 7259 -9881 7981 -9880
rect 6840 -9948 6936 -9932
rect 8252 -9932 8268 -9108
rect 8332 -9932 8348 -9108
rect 9664 -9108 9760 -9092
rect 8671 -9160 9393 -9159
rect 8671 -9880 8672 -9160
rect 9392 -9880 9393 -9160
rect 8671 -9881 9393 -9880
rect 8252 -9948 8348 -9932
rect 9664 -9932 9680 -9108
rect 9744 -9932 9760 -9108
rect 11076 -9108 11172 -9092
rect 10083 -9160 10805 -9159
rect 10083 -9880 10084 -9160
rect 10804 -9880 10805 -9160
rect 10083 -9881 10805 -9880
rect 9664 -9948 9760 -9932
rect 11076 -9932 11092 -9108
rect 11156 -9932 11172 -9108
rect 12488 -9108 12584 -9092
rect 11495 -9160 12217 -9159
rect 11495 -9880 11496 -9160
rect 12216 -9880 12217 -9160
rect 11495 -9881 12217 -9880
rect 11076 -9948 11172 -9932
rect 12488 -9932 12504 -9108
rect 12568 -9932 12584 -9108
rect 13900 -9108 13996 -9092
rect 12907 -9160 13629 -9159
rect 12907 -9880 12908 -9160
rect 13628 -9880 13629 -9160
rect 12907 -9881 13629 -9880
rect 12488 -9948 12584 -9932
rect 13900 -9932 13916 -9108
rect 13980 -9932 13996 -9108
rect 15312 -9108 15408 -9092
rect 14319 -9160 15041 -9159
rect 14319 -9880 14320 -9160
rect 15040 -9880 15041 -9160
rect 14319 -9881 15041 -9880
rect 13900 -9948 13996 -9932
rect 15312 -9932 15328 -9108
rect 15392 -9932 15408 -9108
rect 16724 -9108 16820 -9092
rect 15731 -9160 16453 -9159
rect 15731 -9880 15732 -9160
rect 16452 -9880 16453 -9160
rect 15731 -9881 16453 -9880
rect 15312 -9948 15408 -9932
rect 16724 -9932 16740 -9108
rect 16804 -9932 16820 -9108
rect 18136 -9108 18232 -9092
rect 17143 -9160 17865 -9159
rect 17143 -9880 17144 -9160
rect 17864 -9880 17865 -9160
rect 17143 -9881 17865 -9880
rect 16724 -9948 16820 -9932
rect 18136 -9932 18152 -9108
rect 18216 -9932 18232 -9108
rect 19548 -9108 19644 -9092
rect 18555 -9160 19277 -9159
rect 18555 -9880 18556 -9160
rect 19276 -9880 19277 -9160
rect 18555 -9881 19277 -9880
rect 18136 -9948 18232 -9932
rect 19548 -9932 19564 -9108
rect 19628 -9932 19644 -9108
rect 20960 -9108 21056 -9092
rect 19967 -9160 20689 -9159
rect 19967 -9880 19968 -9160
rect 20688 -9880 20689 -9160
rect 19967 -9881 20689 -9880
rect 19548 -9948 19644 -9932
rect 20960 -9932 20976 -9108
rect 21040 -9932 21056 -9108
rect 22372 -9108 22468 -9092
rect 21379 -9160 22101 -9159
rect 21379 -9880 21380 -9160
rect 22100 -9880 22101 -9160
rect 21379 -9881 22101 -9880
rect 20960 -9948 21056 -9932
rect 22372 -9932 22388 -9108
rect 22452 -9932 22468 -9108
rect 23784 -9108 23880 -9092
rect 22791 -9160 23513 -9159
rect 22791 -9880 22792 -9160
rect 23512 -9880 23513 -9160
rect 22791 -9881 23513 -9880
rect 22372 -9948 22468 -9932
rect 23784 -9932 23800 -9108
rect 23864 -9932 23880 -9108
rect 23784 -9948 23880 -9932
rect -22812 -10228 -22716 -10212
rect -23805 -10280 -23083 -10279
rect -23805 -11000 -23804 -10280
rect -23084 -11000 -23083 -10280
rect -23805 -11001 -23083 -11000
rect -22812 -11052 -22796 -10228
rect -22732 -11052 -22716 -10228
rect -21400 -10228 -21304 -10212
rect -22393 -10280 -21671 -10279
rect -22393 -11000 -22392 -10280
rect -21672 -11000 -21671 -10280
rect -22393 -11001 -21671 -11000
rect -22812 -11068 -22716 -11052
rect -21400 -11052 -21384 -10228
rect -21320 -11052 -21304 -10228
rect -19988 -10228 -19892 -10212
rect -20981 -10280 -20259 -10279
rect -20981 -11000 -20980 -10280
rect -20260 -11000 -20259 -10280
rect -20981 -11001 -20259 -11000
rect -21400 -11068 -21304 -11052
rect -19988 -11052 -19972 -10228
rect -19908 -11052 -19892 -10228
rect -18576 -10228 -18480 -10212
rect -19569 -10280 -18847 -10279
rect -19569 -11000 -19568 -10280
rect -18848 -11000 -18847 -10280
rect -19569 -11001 -18847 -11000
rect -19988 -11068 -19892 -11052
rect -18576 -11052 -18560 -10228
rect -18496 -11052 -18480 -10228
rect -17164 -10228 -17068 -10212
rect -18157 -10280 -17435 -10279
rect -18157 -11000 -18156 -10280
rect -17436 -11000 -17435 -10280
rect -18157 -11001 -17435 -11000
rect -18576 -11068 -18480 -11052
rect -17164 -11052 -17148 -10228
rect -17084 -11052 -17068 -10228
rect -15752 -10228 -15656 -10212
rect -16745 -10280 -16023 -10279
rect -16745 -11000 -16744 -10280
rect -16024 -11000 -16023 -10280
rect -16745 -11001 -16023 -11000
rect -17164 -11068 -17068 -11052
rect -15752 -11052 -15736 -10228
rect -15672 -11052 -15656 -10228
rect -14340 -10228 -14244 -10212
rect -15333 -10280 -14611 -10279
rect -15333 -11000 -15332 -10280
rect -14612 -11000 -14611 -10280
rect -15333 -11001 -14611 -11000
rect -15752 -11068 -15656 -11052
rect -14340 -11052 -14324 -10228
rect -14260 -11052 -14244 -10228
rect -12928 -10228 -12832 -10212
rect -13921 -10280 -13199 -10279
rect -13921 -11000 -13920 -10280
rect -13200 -11000 -13199 -10280
rect -13921 -11001 -13199 -11000
rect -14340 -11068 -14244 -11052
rect -12928 -11052 -12912 -10228
rect -12848 -11052 -12832 -10228
rect -11516 -10228 -11420 -10212
rect -12509 -10280 -11787 -10279
rect -12509 -11000 -12508 -10280
rect -11788 -11000 -11787 -10280
rect -12509 -11001 -11787 -11000
rect -12928 -11068 -12832 -11052
rect -11516 -11052 -11500 -10228
rect -11436 -11052 -11420 -10228
rect -10104 -10228 -10008 -10212
rect -11097 -10280 -10375 -10279
rect -11097 -11000 -11096 -10280
rect -10376 -11000 -10375 -10280
rect -11097 -11001 -10375 -11000
rect -11516 -11068 -11420 -11052
rect -10104 -11052 -10088 -10228
rect -10024 -11052 -10008 -10228
rect -8692 -10228 -8596 -10212
rect -9685 -10280 -8963 -10279
rect -9685 -11000 -9684 -10280
rect -8964 -11000 -8963 -10280
rect -9685 -11001 -8963 -11000
rect -10104 -11068 -10008 -11052
rect -8692 -11052 -8676 -10228
rect -8612 -11052 -8596 -10228
rect -7280 -10228 -7184 -10212
rect -8273 -10280 -7551 -10279
rect -8273 -11000 -8272 -10280
rect -7552 -11000 -7551 -10280
rect -8273 -11001 -7551 -11000
rect -8692 -11068 -8596 -11052
rect -7280 -11052 -7264 -10228
rect -7200 -11052 -7184 -10228
rect -5868 -10228 -5772 -10212
rect -6861 -10280 -6139 -10279
rect -6861 -11000 -6860 -10280
rect -6140 -11000 -6139 -10280
rect -6861 -11001 -6139 -11000
rect -7280 -11068 -7184 -11052
rect -5868 -11052 -5852 -10228
rect -5788 -11052 -5772 -10228
rect -4456 -10228 -4360 -10212
rect -5449 -10280 -4727 -10279
rect -5449 -11000 -5448 -10280
rect -4728 -11000 -4727 -10280
rect -5449 -11001 -4727 -11000
rect -5868 -11068 -5772 -11052
rect -4456 -11052 -4440 -10228
rect -4376 -11052 -4360 -10228
rect -3044 -10228 -2948 -10212
rect -4037 -10280 -3315 -10279
rect -4037 -11000 -4036 -10280
rect -3316 -11000 -3315 -10280
rect -4037 -11001 -3315 -11000
rect -4456 -11068 -4360 -11052
rect -3044 -11052 -3028 -10228
rect -2964 -11052 -2948 -10228
rect -1632 -10228 -1536 -10212
rect -2625 -10280 -1903 -10279
rect -2625 -11000 -2624 -10280
rect -1904 -11000 -1903 -10280
rect -2625 -11001 -1903 -11000
rect -3044 -11068 -2948 -11052
rect -1632 -11052 -1616 -10228
rect -1552 -11052 -1536 -10228
rect -220 -10228 -124 -10212
rect -1213 -10280 -491 -10279
rect -1213 -11000 -1212 -10280
rect -492 -11000 -491 -10280
rect -1213 -11001 -491 -11000
rect -1632 -11068 -1536 -11052
rect -220 -11052 -204 -10228
rect -140 -11052 -124 -10228
rect 1192 -10228 1288 -10212
rect 199 -10280 921 -10279
rect 199 -11000 200 -10280
rect 920 -11000 921 -10280
rect 199 -11001 921 -11000
rect -220 -11068 -124 -11052
rect 1192 -11052 1208 -10228
rect 1272 -11052 1288 -10228
rect 2604 -10228 2700 -10212
rect 1611 -10280 2333 -10279
rect 1611 -11000 1612 -10280
rect 2332 -11000 2333 -10280
rect 1611 -11001 2333 -11000
rect 1192 -11068 1288 -11052
rect 2604 -11052 2620 -10228
rect 2684 -11052 2700 -10228
rect 4016 -10228 4112 -10212
rect 3023 -10280 3745 -10279
rect 3023 -11000 3024 -10280
rect 3744 -11000 3745 -10280
rect 3023 -11001 3745 -11000
rect 2604 -11068 2700 -11052
rect 4016 -11052 4032 -10228
rect 4096 -11052 4112 -10228
rect 5428 -10228 5524 -10212
rect 4435 -10280 5157 -10279
rect 4435 -11000 4436 -10280
rect 5156 -11000 5157 -10280
rect 4435 -11001 5157 -11000
rect 4016 -11068 4112 -11052
rect 5428 -11052 5444 -10228
rect 5508 -11052 5524 -10228
rect 6840 -10228 6936 -10212
rect 5847 -10280 6569 -10279
rect 5847 -11000 5848 -10280
rect 6568 -11000 6569 -10280
rect 5847 -11001 6569 -11000
rect 5428 -11068 5524 -11052
rect 6840 -11052 6856 -10228
rect 6920 -11052 6936 -10228
rect 8252 -10228 8348 -10212
rect 7259 -10280 7981 -10279
rect 7259 -11000 7260 -10280
rect 7980 -11000 7981 -10280
rect 7259 -11001 7981 -11000
rect 6840 -11068 6936 -11052
rect 8252 -11052 8268 -10228
rect 8332 -11052 8348 -10228
rect 9664 -10228 9760 -10212
rect 8671 -10280 9393 -10279
rect 8671 -11000 8672 -10280
rect 9392 -11000 9393 -10280
rect 8671 -11001 9393 -11000
rect 8252 -11068 8348 -11052
rect 9664 -11052 9680 -10228
rect 9744 -11052 9760 -10228
rect 11076 -10228 11172 -10212
rect 10083 -10280 10805 -10279
rect 10083 -11000 10084 -10280
rect 10804 -11000 10805 -10280
rect 10083 -11001 10805 -11000
rect 9664 -11068 9760 -11052
rect 11076 -11052 11092 -10228
rect 11156 -11052 11172 -10228
rect 12488 -10228 12584 -10212
rect 11495 -10280 12217 -10279
rect 11495 -11000 11496 -10280
rect 12216 -11000 12217 -10280
rect 11495 -11001 12217 -11000
rect 11076 -11068 11172 -11052
rect 12488 -11052 12504 -10228
rect 12568 -11052 12584 -10228
rect 13900 -10228 13996 -10212
rect 12907 -10280 13629 -10279
rect 12907 -11000 12908 -10280
rect 13628 -11000 13629 -10280
rect 12907 -11001 13629 -11000
rect 12488 -11068 12584 -11052
rect 13900 -11052 13916 -10228
rect 13980 -11052 13996 -10228
rect 15312 -10228 15408 -10212
rect 14319 -10280 15041 -10279
rect 14319 -11000 14320 -10280
rect 15040 -11000 15041 -10280
rect 14319 -11001 15041 -11000
rect 13900 -11068 13996 -11052
rect 15312 -11052 15328 -10228
rect 15392 -11052 15408 -10228
rect 16724 -10228 16820 -10212
rect 15731 -10280 16453 -10279
rect 15731 -11000 15732 -10280
rect 16452 -11000 16453 -10280
rect 15731 -11001 16453 -11000
rect 15312 -11068 15408 -11052
rect 16724 -11052 16740 -10228
rect 16804 -11052 16820 -10228
rect 18136 -10228 18232 -10212
rect 17143 -10280 17865 -10279
rect 17143 -11000 17144 -10280
rect 17864 -11000 17865 -10280
rect 17143 -11001 17865 -11000
rect 16724 -11068 16820 -11052
rect 18136 -11052 18152 -10228
rect 18216 -11052 18232 -10228
rect 19548 -10228 19644 -10212
rect 18555 -10280 19277 -10279
rect 18555 -11000 18556 -10280
rect 19276 -11000 19277 -10280
rect 18555 -11001 19277 -11000
rect 18136 -11068 18232 -11052
rect 19548 -11052 19564 -10228
rect 19628 -11052 19644 -10228
rect 20960 -10228 21056 -10212
rect 19967 -10280 20689 -10279
rect 19967 -11000 19968 -10280
rect 20688 -11000 20689 -10280
rect 19967 -11001 20689 -11000
rect 19548 -11068 19644 -11052
rect 20960 -11052 20976 -10228
rect 21040 -11052 21056 -10228
rect 22372 -10228 22468 -10212
rect 21379 -10280 22101 -10279
rect 21379 -11000 21380 -10280
rect 22100 -11000 22101 -10280
rect 21379 -11001 22101 -11000
rect 20960 -11068 21056 -11052
rect 22372 -11052 22388 -10228
rect 22452 -11052 22468 -10228
rect 23784 -10228 23880 -10212
rect 22791 -10280 23513 -10279
rect 22791 -11000 22792 -10280
rect 23512 -11000 23513 -10280
rect 22791 -11001 23513 -11000
rect 22372 -11068 22468 -11052
rect 23784 -11052 23800 -10228
rect 23864 -11052 23880 -10228
rect 23784 -11068 23880 -11052
rect -22812 -11348 -22716 -11332
rect -23805 -11400 -23083 -11399
rect -23805 -12120 -23804 -11400
rect -23084 -12120 -23083 -11400
rect -23805 -12121 -23083 -12120
rect -22812 -12172 -22796 -11348
rect -22732 -12172 -22716 -11348
rect -21400 -11348 -21304 -11332
rect -22393 -11400 -21671 -11399
rect -22393 -12120 -22392 -11400
rect -21672 -12120 -21671 -11400
rect -22393 -12121 -21671 -12120
rect -22812 -12188 -22716 -12172
rect -21400 -12172 -21384 -11348
rect -21320 -12172 -21304 -11348
rect -19988 -11348 -19892 -11332
rect -20981 -11400 -20259 -11399
rect -20981 -12120 -20980 -11400
rect -20260 -12120 -20259 -11400
rect -20981 -12121 -20259 -12120
rect -21400 -12188 -21304 -12172
rect -19988 -12172 -19972 -11348
rect -19908 -12172 -19892 -11348
rect -18576 -11348 -18480 -11332
rect -19569 -11400 -18847 -11399
rect -19569 -12120 -19568 -11400
rect -18848 -12120 -18847 -11400
rect -19569 -12121 -18847 -12120
rect -19988 -12188 -19892 -12172
rect -18576 -12172 -18560 -11348
rect -18496 -12172 -18480 -11348
rect -17164 -11348 -17068 -11332
rect -18157 -11400 -17435 -11399
rect -18157 -12120 -18156 -11400
rect -17436 -12120 -17435 -11400
rect -18157 -12121 -17435 -12120
rect -18576 -12188 -18480 -12172
rect -17164 -12172 -17148 -11348
rect -17084 -12172 -17068 -11348
rect -15752 -11348 -15656 -11332
rect -16745 -11400 -16023 -11399
rect -16745 -12120 -16744 -11400
rect -16024 -12120 -16023 -11400
rect -16745 -12121 -16023 -12120
rect -17164 -12188 -17068 -12172
rect -15752 -12172 -15736 -11348
rect -15672 -12172 -15656 -11348
rect -14340 -11348 -14244 -11332
rect -15333 -11400 -14611 -11399
rect -15333 -12120 -15332 -11400
rect -14612 -12120 -14611 -11400
rect -15333 -12121 -14611 -12120
rect -15752 -12188 -15656 -12172
rect -14340 -12172 -14324 -11348
rect -14260 -12172 -14244 -11348
rect -12928 -11348 -12832 -11332
rect -13921 -11400 -13199 -11399
rect -13921 -12120 -13920 -11400
rect -13200 -12120 -13199 -11400
rect -13921 -12121 -13199 -12120
rect -14340 -12188 -14244 -12172
rect -12928 -12172 -12912 -11348
rect -12848 -12172 -12832 -11348
rect -11516 -11348 -11420 -11332
rect -12509 -11400 -11787 -11399
rect -12509 -12120 -12508 -11400
rect -11788 -12120 -11787 -11400
rect -12509 -12121 -11787 -12120
rect -12928 -12188 -12832 -12172
rect -11516 -12172 -11500 -11348
rect -11436 -12172 -11420 -11348
rect -10104 -11348 -10008 -11332
rect -11097 -11400 -10375 -11399
rect -11097 -12120 -11096 -11400
rect -10376 -12120 -10375 -11400
rect -11097 -12121 -10375 -12120
rect -11516 -12188 -11420 -12172
rect -10104 -12172 -10088 -11348
rect -10024 -12172 -10008 -11348
rect -8692 -11348 -8596 -11332
rect -9685 -11400 -8963 -11399
rect -9685 -12120 -9684 -11400
rect -8964 -12120 -8963 -11400
rect -9685 -12121 -8963 -12120
rect -10104 -12188 -10008 -12172
rect -8692 -12172 -8676 -11348
rect -8612 -12172 -8596 -11348
rect -7280 -11348 -7184 -11332
rect -8273 -11400 -7551 -11399
rect -8273 -12120 -8272 -11400
rect -7552 -12120 -7551 -11400
rect -8273 -12121 -7551 -12120
rect -8692 -12188 -8596 -12172
rect -7280 -12172 -7264 -11348
rect -7200 -12172 -7184 -11348
rect -5868 -11348 -5772 -11332
rect -6861 -11400 -6139 -11399
rect -6861 -12120 -6860 -11400
rect -6140 -12120 -6139 -11400
rect -6861 -12121 -6139 -12120
rect -7280 -12188 -7184 -12172
rect -5868 -12172 -5852 -11348
rect -5788 -12172 -5772 -11348
rect -4456 -11348 -4360 -11332
rect -5449 -11400 -4727 -11399
rect -5449 -12120 -5448 -11400
rect -4728 -12120 -4727 -11400
rect -5449 -12121 -4727 -12120
rect -5868 -12188 -5772 -12172
rect -4456 -12172 -4440 -11348
rect -4376 -12172 -4360 -11348
rect -3044 -11348 -2948 -11332
rect -4037 -11400 -3315 -11399
rect -4037 -12120 -4036 -11400
rect -3316 -12120 -3315 -11400
rect -4037 -12121 -3315 -12120
rect -4456 -12188 -4360 -12172
rect -3044 -12172 -3028 -11348
rect -2964 -12172 -2948 -11348
rect -1632 -11348 -1536 -11332
rect -2625 -11400 -1903 -11399
rect -2625 -12120 -2624 -11400
rect -1904 -12120 -1903 -11400
rect -2625 -12121 -1903 -12120
rect -3044 -12188 -2948 -12172
rect -1632 -12172 -1616 -11348
rect -1552 -12172 -1536 -11348
rect -220 -11348 -124 -11332
rect -1213 -11400 -491 -11399
rect -1213 -12120 -1212 -11400
rect -492 -12120 -491 -11400
rect -1213 -12121 -491 -12120
rect -1632 -12188 -1536 -12172
rect -220 -12172 -204 -11348
rect -140 -12172 -124 -11348
rect 1192 -11348 1288 -11332
rect 199 -11400 921 -11399
rect 199 -12120 200 -11400
rect 920 -12120 921 -11400
rect 199 -12121 921 -12120
rect -220 -12188 -124 -12172
rect 1192 -12172 1208 -11348
rect 1272 -12172 1288 -11348
rect 2604 -11348 2700 -11332
rect 1611 -11400 2333 -11399
rect 1611 -12120 1612 -11400
rect 2332 -12120 2333 -11400
rect 1611 -12121 2333 -12120
rect 1192 -12188 1288 -12172
rect 2604 -12172 2620 -11348
rect 2684 -12172 2700 -11348
rect 4016 -11348 4112 -11332
rect 3023 -11400 3745 -11399
rect 3023 -12120 3024 -11400
rect 3744 -12120 3745 -11400
rect 3023 -12121 3745 -12120
rect 2604 -12188 2700 -12172
rect 4016 -12172 4032 -11348
rect 4096 -12172 4112 -11348
rect 5428 -11348 5524 -11332
rect 4435 -11400 5157 -11399
rect 4435 -12120 4436 -11400
rect 5156 -12120 5157 -11400
rect 4435 -12121 5157 -12120
rect 4016 -12188 4112 -12172
rect 5428 -12172 5444 -11348
rect 5508 -12172 5524 -11348
rect 6840 -11348 6936 -11332
rect 5847 -11400 6569 -11399
rect 5847 -12120 5848 -11400
rect 6568 -12120 6569 -11400
rect 5847 -12121 6569 -12120
rect 5428 -12188 5524 -12172
rect 6840 -12172 6856 -11348
rect 6920 -12172 6936 -11348
rect 8252 -11348 8348 -11332
rect 7259 -11400 7981 -11399
rect 7259 -12120 7260 -11400
rect 7980 -12120 7981 -11400
rect 7259 -12121 7981 -12120
rect 6840 -12188 6936 -12172
rect 8252 -12172 8268 -11348
rect 8332 -12172 8348 -11348
rect 9664 -11348 9760 -11332
rect 8671 -11400 9393 -11399
rect 8671 -12120 8672 -11400
rect 9392 -12120 9393 -11400
rect 8671 -12121 9393 -12120
rect 8252 -12188 8348 -12172
rect 9664 -12172 9680 -11348
rect 9744 -12172 9760 -11348
rect 11076 -11348 11172 -11332
rect 10083 -11400 10805 -11399
rect 10083 -12120 10084 -11400
rect 10804 -12120 10805 -11400
rect 10083 -12121 10805 -12120
rect 9664 -12188 9760 -12172
rect 11076 -12172 11092 -11348
rect 11156 -12172 11172 -11348
rect 12488 -11348 12584 -11332
rect 11495 -11400 12217 -11399
rect 11495 -12120 11496 -11400
rect 12216 -12120 12217 -11400
rect 11495 -12121 12217 -12120
rect 11076 -12188 11172 -12172
rect 12488 -12172 12504 -11348
rect 12568 -12172 12584 -11348
rect 13900 -11348 13996 -11332
rect 12907 -11400 13629 -11399
rect 12907 -12120 12908 -11400
rect 13628 -12120 13629 -11400
rect 12907 -12121 13629 -12120
rect 12488 -12188 12584 -12172
rect 13900 -12172 13916 -11348
rect 13980 -12172 13996 -11348
rect 15312 -11348 15408 -11332
rect 14319 -11400 15041 -11399
rect 14319 -12120 14320 -11400
rect 15040 -12120 15041 -11400
rect 14319 -12121 15041 -12120
rect 13900 -12188 13996 -12172
rect 15312 -12172 15328 -11348
rect 15392 -12172 15408 -11348
rect 16724 -11348 16820 -11332
rect 15731 -11400 16453 -11399
rect 15731 -12120 15732 -11400
rect 16452 -12120 16453 -11400
rect 15731 -12121 16453 -12120
rect 15312 -12188 15408 -12172
rect 16724 -12172 16740 -11348
rect 16804 -12172 16820 -11348
rect 18136 -11348 18232 -11332
rect 17143 -11400 17865 -11399
rect 17143 -12120 17144 -11400
rect 17864 -12120 17865 -11400
rect 17143 -12121 17865 -12120
rect 16724 -12188 16820 -12172
rect 18136 -12172 18152 -11348
rect 18216 -12172 18232 -11348
rect 19548 -11348 19644 -11332
rect 18555 -11400 19277 -11399
rect 18555 -12120 18556 -11400
rect 19276 -12120 19277 -11400
rect 18555 -12121 19277 -12120
rect 18136 -12188 18232 -12172
rect 19548 -12172 19564 -11348
rect 19628 -12172 19644 -11348
rect 20960 -11348 21056 -11332
rect 19967 -11400 20689 -11399
rect 19967 -12120 19968 -11400
rect 20688 -12120 20689 -11400
rect 19967 -12121 20689 -12120
rect 19548 -12188 19644 -12172
rect 20960 -12172 20976 -11348
rect 21040 -12172 21056 -11348
rect 22372 -11348 22468 -11332
rect 21379 -11400 22101 -11399
rect 21379 -12120 21380 -11400
rect 22100 -12120 22101 -11400
rect 21379 -12121 22101 -12120
rect 20960 -12188 21056 -12172
rect 22372 -12172 22388 -11348
rect 22452 -12172 22468 -11348
rect 23784 -11348 23880 -11332
rect 22791 -11400 23513 -11399
rect 22791 -12120 22792 -11400
rect 23512 -12120 23513 -11400
rect 22791 -12121 23513 -12120
rect 22372 -12188 22468 -12172
rect 23784 -12172 23800 -11348
rect 23864 -12172 23880 -11348
rect 23784 -12188 23880 -12172
rect -22812 -12468 -22716 -12452
rect -23805 -12520 -23083 -12519
rect -23805 -13240 -23804 -12520
rect -23084 -13240 -23083 -12520
rect -23805 -13241 -23083 -13240
rect -22812 -13292 -22796 -12468
rect -22732 -13292 -22716 -12468
rect -21400 -12468 -21304 -12452
rect -22393 -12520 -21671 -12519
rect -22393 -13240 -22392 -12520
rect -21672 -13240 -21671 -12520
rect -22393 -13241 -21671 -13240
rect -22812 -13308 -22716 -13292
rect -21400 -13292 -21384 -12468
rect -21320 -13292 -21304 -12468
rect -19988 -12468 -19892 -12452
rect -20981 -12520 -20259 -12519
rect -20981 -13240 -20980 -12520
rect -20260 -13240 -20259 -12520
rect -20981 -13241 -20259 -13240
rect -21400 -13308 -21304 -13292
rect -19988 -13292 -19972 -12468
rect -19908 -13292 -19892 -12468
rect -18576 -12468 -18480 -12452
rect -19569 -12520 -18847 -12519
rect -19569 -13240 -19568 -12520
rect -18848 -13240 -18847 -12520
rect -19569 -13241 -18847 -13240
rect -19988 -13308 -19892 -13292
rect -18576 -13292 -18560 -12468
rect -18496 -13292 -18480 -12468
rect -17164 -12468 -17068 -12452
rect -18157 -12520 -17435 -12519
rect -18157 -13240 -18156 -12520
rect -17436 -13240 -17435 -12520
rect -18157 -13241 -17435 -13240
rect -18576 -13308 -18480 -13292
rect -17164 -13292 -17148 -12468
rect -17084 -13292 -17068 -12468
rect -15752 -12468 -15656 -12452
rect -16745 -12520 -16023 -12519
rect -16745 -13240 -16744 -12520
rect -16024 -13240 -16023 -12520
rect -16745 -13241 -16023 -13240
rect -17164 -13308 -17068 -13292
rect -15752 -13292 -15736 -12468
rect -15672 -13292 -15656 -12468
rect -14340 -12468 -14244 -12452
rect -15333 -12520 -14611 -12519
rect -15333 -13240 -15332 -12520
rect -14612 -13240 -14611 -12520
rect -15333 -13241 -14611 -13240
rect -15752 -13308 -15656 -13292
rect -14340 -13292 -14324 -12468
rect -14260 -13292 -14244 -12468
rect -12928 -12468 -12832 -12452
rect -13921 -12520 -13199 -12519
rect -13921 -13240 -13920 -12520
rect -13200 -13240 -13199 -12520
rect -13921 -13241 -13199 -13240
rect -14340 -13308 -14244 -13292
rect -12928 -13292 -12912 -12468
rect -12848 -13292 -12832 -12468
rect -11516 -12468 -11420 -12452
rect -12509 -12520 -11787 -12519
rect -12509 -13240 -12508 -12520
rect -11788 -13240 -11787 -12520
rect -12509 -13241 -11787 -13240
rect -12928 -13308 -12832 -13292
rect -11516 -13292 -11500 -12468
rect -11436 -13292 -11420 -12468
rect -10104 -12468 -10008 -12452
rect -11097 -12520 -10375 -12519
rect -11097 -13240 -11096 -12520
rect -10376 -13240 -10375 -12520
rect -11097 -13241 -10375 -13240
rect -11516 -13308 -11420 -13292
rect -10104 -13292 -10088 -12468
rect -10024 -13292 -10008 -12468
rect -8692 -12468 -8596 -12452
rect -9685 -12520 -8963 -12519
rect -9685 -13240 -9684 -12520
rect -8964 -13240 -8963 -12520
rect -9685 -13241 -8963 -13240
rect -10104 -13308 -10008 -13292
rect -8692 -13292 -8676 -12468
rect -8612 -13292 -8596 -12468
rect -7280 -12468 -7184 -12452
rect -8273 -12520 -7551 -12519
rect -8273 -13240 -8272 -12520
rect -7552 -13240 -7551 -12520
rect -8273 -13241 -7551 -13240
rect -8692 -13308 -8596 -13292
rect -7280 -13292 -7264 -12468
rect -7200 -13292 -7184 -12468
rect -5868 -12468 -5772 -12452
rect -6861 -12520 -6139 -12519
rect -6861 -13240 -6860 -12520
rect -6140 -13240 -6139 -12520
rect -6861 -13241 -6139 -13240
rect -7280 -13308 -7184 -13292
rect -5868 -13292 -5852 -12468
rect -5788 -13292 -5772 -12468
rect -4456 -12468 -4360 -12452
rect -5449 -12520 -4727 -12519
rect -5449 -13240 -5448 -12520
rect -4728 -13240 -4727 -12520
rect -5449 -13241 -4727 -13240
rect -5868 -13308 -5772 -13292
rect -4456 -13292 -4440 -12468
rect -4376 -13292 -4360 -12468
rect -3044 -12468 -2948 -12452
rect -4037 -12520 -3315 -12519
rect -4037 -13240 -4036 -12520
rect -3316 -13240 -3315 -12520
rect -4037 -13241 -3315 -13240
rect -4456 -13308 -4360 -13292
rect -3044 -13292 -3028 -12468
rect -2964 -13292 -2948 -12468
rect -1632 -12468 -1536 -12452
rect -2625 -12520 -1903 -12519
rect -2625 -13240 -2624 -12520
rect -1904 -13240 -1903 -12520
rect -2625 -13241 -1903 -13240
rect -3044 -13308 -2948 -13292
rect -1632 -13292 -1616 -12468
rect -1552 -13292 -1536 -12468
rect -220 -12468 -124 -12452
rect -1213 -12520 -491 -12519
rect -1213 -13240 -1212 -12520
rect -492 -13240 -491 -12520
rect -1213 -13241 -491 -13240
rect -1632 -13308 -1536 -13292
rect -220 -13292 -204 -12468
rect -140 -13292 -124 -12468
rect 1192 -12468 1288 -12452
rect 199 -12520 921 -12519
rect 199 -13240 200 -12520
rect 920 -13240 921 -12520
rect 199 -13241 921 -13240
rect -220 -13308 -124 -13292
rect 1192 -13292 1208 -12468
rect 1272 -13292 1288 -12468
rect 2604 -12468 2700 -12452
rect 1611 -12520 2333 -12519
rect 1611 -13240 1612 -12520
rect 2332 -13240 2333 -12520
rect 1611 -13241 2333 -13240
rect 1192 -13308 1288 -13292
rect 2604 -13292 2620 -12468
rect 2684 -13292 2700 -12468
rect 4016 -12468 4112 -12452
rect 3023 -12520 3745 -12519
rect 3023 -13240 3024 -12520
rect 3744 -13240 3745 -12520
rect 3023 -13241 3745 -13240
rect 2604 -13308 2700 -13292
rect 4016 -13292 4032 -12468
rect 4096 -13292 4112 -12468
rect 5428 -12468 5524 -12452
rect 4435 -12520 5157 -12519
rect 4435 -13240 4436 -12520
rect 5156 -13240 5157 -12520
rect 4435 -13241 5157 -13240
rect 4016 -13308 4112 -13292
rect 5428 -13292 5444 -12468
rect 5508 -13292 5524 -12468
rect 6840 -12468 6936 -12452
rect 5847 -12520 6569 -12519
rect 5847 -13240 5848 -12520
rect 6568 -13240 6569 -12520
rect 5847 -13241 6569 -13240
rect 5428 -13308 5524 -13292
rect 6840 -13292 6856 -12468
rect 6920 -13292 6936 -12468
rect 8252 -12468 8348 -12452
rect 7259 -12520 7981 -12519
rect 7259 -13240 7260 -12520
rect 7980 -13240 7981 -12520
rect 7259 -13241 7981 -13240
rect 6840 -13308 6936 -13292
rect 8252 -13292 8268 -12468
rect 8332 -13292 8348 -12468
rect 9664 -12468 9760 -12452
rect 8671 -12520 9393 -12519
rect 8671 -13240 8672 -12520
rect 9392 -13240 9393 -12520
rect 8671 -13241 9393 -13240
rect 8252 -13308 8348 -13292
rect 9664 -13292 9680 -12468
rect 9744 -13292 9760 -12468
rect 11076 -12468 11172 -12452
rect 10083 -12520 10805 -12519
rect 10083 -13240 10084 -12520
rect 10804 -13240 10805 -12520
rect 10083 -13241 10805 -13240
rect 9664 -13308 9760 -13292
rect 11076 -13292 11092 -12468
rect 11156 -13292 11172 -12468
rect 12488 -12468 12584 -12452
rect 11495 -12520 12217 -12519
rect 11495 -13240 11496 -12520
rect 12216 -13240 12217 -12520
rect 11495 -13241 12217 -13240
rect 11076 -13308 11172 -13292
rect 12488 -13292 12504 -12468
rect 12568 -13292 12584 -12468
rect 13900 -12468 13996 -12452
rect 12907 -12520 13629 -12519
rect 12907 -13240 12908 -12520
rect 13628 -13240 13629 -12520
rect 12907 -13241 13629 -13240
rect 12488 -13308 12584 -13292
rect 13900 -13292 13916 -12468
rect 13980 -13292 13996 -12468
rect 15312 -12468 15408 -12452
rect 14319 -12520 15041 -12519
rect 14319 -13240 14320 -12520
rect 15040 -13240 15041 -12520
rect 14319 -13241 15041 -13240
rect 13900 -13308 13996 -13292
rect 15312 -13292 15328 -12468
rect 15392 -13292 15408 -12468
rect 16724 -12468 16820 -12452
rect 15731 -12520 16453 -12519
rect 15731 -13240 15732 -12520
rect 16452 -13240 16453 -12520
rect 15731 -13241 16453 -13240
rect 15312 -13308 15408 -13292
rect 16724 -13292 16740 -12468
rect 16804 -13292 16820 -12468
rect 18136 -12468 18232 -12452
rect 17143 -12520 17865 -12519
rect 17143 -13240 17144 -12520
rect 17864 -13240 17865 -12520
rect 17143 -13241 17865 -13240
rect 16724 -13308 16820 -13292
rect 18136 -13292 18152 -12468
rect 18216 -13292 18232 -12468
rect 19548 -12468 19644 -12452
rect 18555 -12520 19277 -12519
rect 18555 -13240 18556 -12520
rect 19276 -13240 19277 -12520
rect 18555 -13241 19277 -13240
rect 18136 -13308 18232 -13292
rect 19548 -13292 19564 -12468
rect 19628 -13292 19644 -12468
rect 20960 -12468 21056 -12452
rect 19967 -12520 20689 -12519
rect 19967 -13240 19968 -12520
rect 20688 -13240 20689 -12520
rect 19967 -13241 20689 -13240
rect 19548 -13308 19644 -13292
rect 20960 -13292 20976 -12468
rect 21040 -13292 21056 -12468
rect 22372 -12468 22468 -12452
rect 21379 -12520 22101 -12519
rect 21379 -13240 21380 -12520
rect 22100 -13240 22101 -12520
rect 21379 -13241 22101 -13240
rect 20960 -13308 21056 -13292
rect 22372 -13292 22388 -12468
rect 22452 -13292 22468 -12468
rect 23784 -12468 23880 -12452
rect 22791 -12520 23513 -12519
rect 22791 -13240 22792 -12520
rect 23512 -13240 23513 -12520
rect 22791 -13241 23513 -13240
rect 22372 -13308 22468 -13292
rect 23784 -13292 23800 -12468
rect 23864 -13292 23880 -12468
rect 23784 -13308 23880 -13292
rect -22812 -13588 -22716 -13572
rect -23805 -13640 -23083 -13639
rect -23805 -14360 -23804 -13640
rect -23084 -14360 -23083 -13640
rect -23805 -14361 -23083 -14360
rect -22812 -14412 -22796 -13588
rect -22732 -14412 -22716 -13588
rect -21400 -13588 -21304 -13572
rect -22393 -13640 -21671 -13639
rect -22393 -14360 -22392 -13640
rect -21672 -14360 -21671 -13640
rect -22393 -14361 -21671 -14360
rect -22812 -14428 -22716 -14412
rect -21400 -14412 -21384 -13588
rect -21320 -14412 -21304 -13588
rect -19988 -13588 -19892 -13572
rect -20981 -13640 -20259 -13639
rect -20981 -14360 -20980 -13640
rect -20260 -14360 -20259 -13640
rect -20981 -14361 -20259 -14360
rect -21400 -14428 -21304 -14412
rect -19988 -14412 -19972 -13588
rect -19908 -14412 -19892 -13588
rect -18576 -13588 -18480 -13572
rect -19569 -13640 -18847 -13639
rect -19569 -14360 -19568 -13640
rect -18848 -14360 -18847 -13640
rect -19569 -14361 -18847 -14360
rect -19988 -14428 -19892 -14412
rect -18576 -14412 -18560 -13588
rect -18496 -14412 -18480 -13588
rect -17164 -13588 -17068 -13572
rect -18157 -13640 -17435 -13639
rect -18157 -14360 -18156 -13640
rect -17436 -14360 -17435 -13640
rect -18157 -14361 -17435 -14360
rect -18576 -14428 -18480 -14412
rect -17164 -14412 -17148 -13588
rect -17084 -14412 -17068 -13588
rect -15752 -13588 -15656 -13572
rect -16745 -13640 -16023 -13639
rect -16745 -14360 -16744 -13640
rect -16024 -14360 -16023 -13640
rect -16745 -14361 -16023 -14360
rect -17164 -14428 -17068 -14412
rect -15752 -14412 -15736 -13588
rect -15672 -14412 -15656 -13588
rect -14340 -13588 -14244 -13572
rect -15333 -13640 -14611 -13639
rect -15333 -14360 -15332 -13640
rect -14612 -14360 -14611 -13640
rect -15333 -14361 -14611 -14360
rect -15752 -14428 -15656 -14412
rect -14340 -14412 -14324 -13588
rect -14260 -14412 -14244 -13588
rect -12928 -13588 -12832 -13572
rect -13921 -13640 -13199 -13639
rect -13921 -14360 -13920 -13640
rect -13200 -14360 -13199 -13640
rect -13921 -14361 -13199 -14360
rect -14340 -14428 -14244 -14412
rect -12928 -14412 -12912 -13588
rect -12848 -14412 -12832 -13588
rect -11516 -13588 -11420 -13572
rect -12509 -13640 -11787 -13639
rect -12509 -14360 -12508 -13640
rect -11788 -14360 -11787 -13640
rect -12509 -14361 -11787 -14360
rect -12928 -14428 -12832 -14412
rect -11516 -14412 -11500 -13588
rect -11436 -14412 -11420 -13588
rect -10104 -13588 -10008 -13572
rect -11097 -13640 -10375 -13639
rect -11097 -14360 -11096 -13640
rect -10376 -14360 -10375 -13640
rect -11097 -14361 -10375 -14360
rect -11516 -14428 -11420 -14412
rect -10104 -14412 -10088 -13588
rect -10024 -14412 -10008 -13588
rect -8692 -13588 -8596 -13572
rect -9685 -13640 -8963 -13639
rect -9685 -14360 -9684 -13640
rect -8964 -14360 -8963 -13640
rect -9685 -14361 -8963 -14360
rect -10104 -14428 -10008 -14412
rect -8692 -14412 -8676 -13588
rect -8612 -14412 -8596 -13588
rect -7280 -13588 -7184 -13572
rect -8273 -13640 -7551 -13639
rect -8273 -14360 -8272 -13640
rect -7552 -14360 -7551 -13640
rect -8273 -14361 -7551 -14360
rect -8692 -14428 -8596 -14412
rect -7280 -14412 -7264 -13588
rect -7200 -14412 -7184 -13588
rect -5868 -13588 -5772 -13572
rect -6861 -13640 -6139 -13639
rect -6861 -14360 -6860 -13640
rect -6140 -14360 -6139 -13640
rect -6861 -14361 -6139 -14360
rect -7280 -14428 -7184 -14412
rect -5868 -14412 -5852 -13588
rect -5788 -14412 -5772 -13588
rect -4456 -13588 -4360 -13572
rect -5449 -13640 -4727 -13639
rect -5449 -14360 -5448 -13640
rect -4728 -14360 -4727 -13640
rect -5449 -14361 -4727 -14360
rect -5868 -14428 -5772 -14412
rect -4456 -14412 -4440 -13588
rect -4376 -14412 -4360 -13588
rect -3044 -13588 -2948 -13572
rect -4037 -13640 -3315 -13639
rect -4037 -14360 -4036 -13640
rect -3316 -14360 -3315 -13640
rect -4037 -14361 -3315 -14360
rect -4456 -14428 -4360 -14412
rect -3044 -14412 -3028 -13588
rect -2964 -14412 -2948 -13588
rect -1632 -13588 -1536 -13572
rect -2625 -13640 -1903 -13639
rect -2625 -14360 -2624 -13640
rect -1904 -14360 -1903 -13640
rect -2625 -14361 -1903 -14360
rect -3044 -14428 -2948 -14412
rect -1632 -14412 -1616 -13588
rect -1552 -14412 -1536 -13588
rect -220 -13588 -124 -13572
rect -1213 -13640 -491 -13639
rect -1213 -14360 -1212 -13640
rect -492 -14360 -491 -13640
rect -1213 -14361 -491 -14360
rect -1632 -14428 -1536 -14412
rect -220 -14412 -204 -13588
rect -140 -14412 -124 -13588
rect 1192 -13588 1288 -13572
rect 199 -13640 921 -13639
rect 199 -14360 200 -13640
rect 920 -14360 921 -13640
rect 199 -14361 921 -14360
rect -220 -14428 -124 -14412
rect 1192 -14412 1208 -13588
rect 1272 -14412 1288 -13588
rect 2604 -13588 2700 -13572
rect 1611 -13640 2333 -13639
rect 1611 -14360 1612 -13640
rect 2332 -14360 2333 -13640
rect 1611 -14361 2333 -14360
rect 1192 -14428 1288 -14412
rect 2604 -14412 2620 -13588
rect 2684 -14412 2700 -13588
rect 4016 -13588 4112 -13572
rect 3023 -13640 3745 -13639
rect 3023 -14360 3024 -13640
rect 3744 -14360 3745 -13640
rect 3023 -14361 3745 -14360
rect 2604 -14428 2700 -14412
rect 4016 -14412 4032 -13588
rect 4096 -14412 4112 -13588
rect 5428 -13588 5524 -13572
rect 4435 -13640 5157 -13639
rect 4435 -14360 4436 -13640
rect 5156 -14360 5157 -13640
rect 4435 -14361 5157 -14360
rect 4016 -14428 4112 -14412
rect 5428 -14412 5444 -13588
rect 5508 -14412 5524 -13588
rect 6840 -13588 6936 -13572
rect 5847 -13640 6569 -13639
rect 5847 -14360 5848 -13640
rect 6568 -14360 6569 -13640
rect 5847 -14361 6569 -14360
rect 5428 -14428 5524 -14412
rect 6840 -14412 6856 -13588
rect 6920 -14412 6936 -13588
rect 8252 -13588 8348 -13572
rect 7259 -13640 7981 -13639
rect 7259 -14360 7260 -13640
rect 7980 -14360 7981 -13640
rect 7259 -14361 7981 -14360
rect 6840 -14428 6936 -14412
rect 8252 -14412 8268 -13588
rect 8332 -14412 8348 -13588
rect 9664 -13588 9760 -13572
rect 8671 -13640 9393 -13639
rect 8671 -14360 8672 -13640
rect 9392 -14360 9393 -13640
rect 8671 -14361 9393 -14360
rect 8252 -14428 8348 -14412
rect 9664 -14412 9680 -13588
rect 9744 -14412 9760 -13588
rect 11076 -13588 11172 -13572
rect 10083 -13640 10805 -13639
rect 10083 -14360 10084 -13640
rect 10804 -14360 10805 -13640
rect 10083 -14361 10805 -14360
rect 9664 -14428 9760 -14412
rect 11076 -14412 11092 -13588
rect 11156 -14412 11172 -13588
rect 12488 -13588 12584 -13572
rect 11495 -13640 12217 -13639
rect 11495 -14360 11496 -13640
rect 12216 -14360 12217 -13640
rect 11495 -14361 12217 -14360
rect 11076 -14428 11172 -14412
rect 12488 -14412 12504 -13588
rect 12568 -14412 12584 -13588
rect 13900 -13588 13996 -13572
rect 12907 -13640 13629 -13639
rect 12907 -14360 12908 -13640
rect 13628 -14360 13629 -13640
rect 12907 -14361 13629 -14360
rect 12488 -14428 12584 -14412
rect 13900 -14412 13916 -13588
rect 13980 -14412 13996 -13588
rect 15312 -13588 15408 -13572
rect 14319 -13640 15041 -13639
rect 14319 -14360 14320 -13640
rect 15040 -14360 15041 -13640
rect 14319 -14361 15041 -14360
rect 13900 -14428 13996 -14412
rect 15312 -14412 15328 -13588
rect 15392 -14412 15408 -13588
rect 16724 -13588 16820 -13572
rect 15731 -13640 16453 -13639
rect 15731 -14360 15732 -13640
rect 16452 -14360 16453 -13640
rect 15731 -14361 16453 -14360
rect 15312 -14428 15408 -14412
rect 16724 -14412 16740 -13588
rect 16804 -14412 16820 -13588
rect 18136 -13588 18232 -13572
rect 17143 -13640 17865 -13639
rect 17143 -14360 17144 -13640
rect 17864 -14360 17865 -13640
rect 17143 -14361 17865 -14360
rect 16724 -14428 16820 -14412
rect 18136 -14412 18152 -13588
rect 18216 -14412 18232 -13588
rect 19548 -13588 19644 -13572
rect 18555 -13640 19277 -13639
rect 18555 -14360 18556 -13640
rect 19276 -14360 19277 -13640
rect 18555 -14361 19277 -14360
rect 18136 -14428 18232 -14412
rect 19548 -14412 19564 -13588
rect 19628 -14412 19644 -13588
rect 20960 -13588 21056 -13572
rect 19967 -13640 20689 -13639
rect 19967 -14360 19968 -13640
rect 20688 -14360 20689 -13640
rect 19967 -14361 20689 -14360
rect 19548 -14428 19644 -14412
rect 20960 -14412 20976 -13588
rect 21040 -14412 21056 -13588
rect 22372 -13588 22468 -13572
rect 21379 -13640 22101 -13639
rect 21379 -14360 21380 -13640
rect 22100 -14360 22101 -13640
rect 21379 -14361 22101 -14360
rect 20960 -14428 21056 -14412
rect 22372 -14412 22388 -13588
rect 22452 -14412 22468 -13588
rect 23784 -13588 23880 -13572
rect 22791 -13640 23513 -13639
rect 22791 -14360 22792 -13640
rect 23512 -14360 23513 -13640
rect 22791 -14361 23513 -14360
rect 22372 -14428 22468 -14412
rect 23784 -14412 23800 -13588
rect 23864 -14412 23880 -13588
rect 23784 -14428 23880 -14412
rect -22812 -14708 -22716 -14692
rect -23805 -14760 -23083 -14759
rect -23805 -15480 -23804 -14760
rect -23084 -15480 -23083 -14760
rect -23805 -15481 -23083 -15480
rect -22812 -15532 -22796 -14708
rect -22732 -15532 -22716 -14708
rect -21400 -14708 -21304 -14692
rect -22393 -14760 -21671 -14759
rect -22393 -15480 -22392 -14760
rect -21672 -15480 -21671 -14760
rect -22393 -15481 -21671 -15480
rect -22812 -15548 -22716 -15532
rect -21400 -15532 -21384 -14708
rect -21320 -15532 -21304 -14708
rect -19988 -14708 -19892 -14692
rect -20981 -14760 -20259 -14759
rect -20981 -15480 -20980 -14760
rect -20260 -15480 -20259 -14760
rect -20981 -15481 -20259 -15480
rect -21400 -15548 -21304 -15532
rect -19988 -15532 -19972 -14708
rect -19908 -15532 -19892 -14708
rect -18576 -14708 -18480 -14692
rect -19569 -14760 -18847 -14759
rect -19569 -15480 -19568 -14760
rect -18848 -15480 -18847 -14760
rect -19569 -15481 -18847 -15480
rect -19988 -15548 -19892 -15532
rect -18576 -15532 -18560 -14708
rect -18496 -15532 -18480 -14708
rect -17164 -14708 -17068 -14692
rect -18157 -14760 -17435 -14759
rect -18157 -15480 -18156 -14760
rect -17436 -15480 -17435 -14760
rect -18157 -15481 -17435 -15480
rect -18576 -15548 -18480 -15532
rect -17164 -15532 -17148 -14708
rect -17084 -15532 -17068 -14708
rect -15752 -14708 -15656 -14692
rect -16745 -14760 -16023 -14759
rect -16745 -15480 -16744 -14760
rect -16024 -15480 -16023 -14760
rect -16745 -15481 -16023 -15480
rect -17164 -15548 -17068 -15532
rect -15752 -15532 -15736 -14708
rect -15672 -15532 -15656 -14708
rect -14340 -14708 -14244 -14692
rect -15333 -14760 -14611 -14759
rect -15333 -15480 -15332 -14760
rect -14612 -15480 -14611 -14760
rect -15333 -15481 -14611 -15480
rect -15752 -15548 -15656 -15532
rect -14340 -15532 -14324 -14708
rect -14260 -15532 -14244 -14708
rect -12928 -14708 -12832 -14692
rect -13921 -14760 -13199 -14759
rect -13921 -15480 -13920 -14760
rect -13200 -15480 -13199 -14760
rect -13921 -15481 -13199 -15480
rect -14340 -15548 -14244 -15532
rect -12928 -15532 -12912 -14708
rect -12848 -15532 -12832 -14708
rect -11516 -14708 -11420 -14692
rect -12509 -14760 -11787 -14759
rect -12509 -15480 -12508 -14760
rect -11788 -15480 -11787 -14760
rect -12509 -15481 -11787 -15480
rect -12928 -15548 -12832 -15532
rect -11516 -15532 -11500 -14708
rect -11436 -15532 -11420 -14708
rect -10104 -14708 -10008 -14692
rect -11097 -14760 -10375 -14759
rect -11097 -15480 -11096 -14760
rect -10376 -15480 -10375 -14760
rect -11097 -15481 -10375 -15480
rect -11516 -15548 -11420 -15532
rect -10104 -15532 -10088 -14708
rect -10024 -15532 -10008 -14708
rect -8692 -14708 -8596 -14692
rect -9685 -14760 -8963 -14759
rect -9685 -15480 -9684 -14760
rect -8964 -15480 -8963 -14760
rect -9685 -15481 -8963 -15480
rect -10104 -15548 -10008 -15532
rect -8692 -15532 -8676 -14708
rect -8612 -15532 -8596 -14708
rect -7280 -14708 -7184 -14692
rect -8273 -14760 -7551 -14759
rect -8273 -15480 -8272 -14760
rect -7552 -15480 -7551 -14760
rect -8273 -15481 -7551 -15480
rect -8692 -15548 -8596 -15532
rect -7280 -15532 -7264 -14708
rect -7200 -15532 -7184 -14708
rect -5868 -14708 -5772 -14692
rect -6861 -14760 -6139 -14759
rect -6861 -15480 -6860 -14760
rect -6140 -15480 -6139 -14760
rect -6861 -15481 -6139 -15480
rect -7280 -15548 -7184 -15532
rect -5868 -15532 -5852 -14708
rect -5788 -15532 -5772 -14708
rect -4456 -14708 -4360 -14692
rect -5449 -14760 -4727 -14759
rect -5449 -15480 -5448 -14760
rect -4728 -15480 -4727 -14760
rect -5449 -15481 -4727 -15480
rect -5868 -15548 -5772 -15532
rect -4456 -15532 -4440 -14708
rect -4376 -15532 -4360 -14708
rect -3044 -14708 -2948 -14692
rect -4037 -14760 -3315 -14759
rect -4037 -15480 -4036 -14760
rect -3316 -15480 -3315 -14760
rect -4037 -15481 -3315 -15480
rect -4456 -15548 -4360 -15532
rect -3044 -15532 -3028 -14708
rect -2964 -15532 -2948 -14708
rect -1632 -14708 -1536 -14692
rect -2625 -14760 -1903 -14759
rect -2625 -15480 -2624 -14760
rect -1904 -15480 -1903 -14760
rect -2625 -15481 -1903 -15480
rect -3044 -15548 -2948 -15532
rect -1632 -15532 -1616 -14708
rect -1552 -15532 -1536 -14708
rect -220 -14708 -124 -14692
rect -1213 -14760 -491 -14759
rect -1213 -15480 -1212 -14760
rect -492 -15480 -491 -14760
rect -1213 -15481 -491 -15480
rect -1632 -15548 -1536 -15532
rect -220 -15532 -204 -14708
rect -140 -15532 -124 -14708
rect 1192 -14708 1288 -14692
rect 199 -14760 921 -14759
rect 199 -15480 200 -14760
rect 920 -15480 921 -14760
rect 199 -15481 921 -15480
rect -220 -15548 -124 -15532
rect 1192 -15532 1208 -14708
rect 1272 -15532 1288 -14708
rect 2604 -14708 2700 -14692
rect 1611 -14760 2333 -14759
rect 1611 -15480 1612 -14760
rect 2332 -15480 2333 -14760
rect 1611 -15481 2333 -15480
rect 1192 -15548 1288 -15532
rect 2604 -15532 2620 -14708
rect 2684 -15532 2700 -14708
rect 4016 -14708 4112 -14692
rect 3023 -14760 3745 -14759
rect 3023 -15480 3024 -14760
rect 3744 -15480 3745 -14760
rect 3023 -15481 3745 -15480
rect 2604 -15548 2700 -15532
rect 4016 -15532 4032 -14708
rect 4096 -15532 4112 -14708
rect 5428 -14708 5524 -14692
rect 4435 -14760 5157 -14759
rect 4435 -15480 4436 -14760
rect 5156 -15480 5157 -14760
rect 4435 -15481 5157 -15480
rect 4016 -15548 4112 -15532
rect 5428 -15532 5444 -14708
rect 5508 -15532 5524 -14708
rect 6840 -14708 6936 -14692
rect 5847 -14760 6569 -14759
rect 5847 -15480 5848 -14760
rect 6568 -15480 6569 -14760
rect 5847 -15481 6569 -15480
rect 5428 -15548 5524 -15532
rect 6840 -15532 6856 -14708
rect 6920 -15532 6936 -14708
rect 8252 -14708 8348 -14692
rect 7259 -14760 7981 -14759
rect 7259 -15480 7260 -14760
rect 7980 -15480 7981 -14760
rect 7259 -15481 7981 -15480
rect 6840 -15548 6936 -15532
rect 8252 -15532 8268 -14708
rect 8332 -15532 8348 -14708
rect 9664 -14708 9760 -14692
rect 8671 -14760 9393 -14759
rect 8671 -15480 8672 -14760
rect 9392 -15480 9393 -14760
rect 8671 -15481 9393 -15480
rect 8252 -15548 8348 -15532
rect 9664 -15532 9680 -14708
rect 9744 -15532 9760 -14708
rect 11076 -14708 11172 -14692
rect 10083 -14760 10805 -14759
rect 10083 -15480 10084 -14760
rect 10804 -15480 10805 -14760
rect 10083 -15481 10805 -15480
rect 9664 -15548 9760 -15532
rect 11076 -15532 11092 -14708
rect 11156 -15532 11172 -14708
rect 12488 -14708 12584 -14692
rect 11495 -14760 12217 -14759
rect 11495 -15480 11496 -14760
rect 12216 -15480 12217 -14760
rect 11495 -15481 12217 -15480
rect 11076 -15548 11172 -15532
rect 12488 -15532 12504 -14708
rect 12568 -15532 12584 -14708
rect 13900 -14708 13996 -14692
rect 12907 -14760 13629 -14759
rect 12907 -15480 12908 -14760
rect 13628 -15480 13629 -14760
rect 12907 -15481 13629 -15480
rect 12488 -15548 12584 -15532
rect 13900 -15532 13916 -14708
rect 13980 -15532 13996 -14708
rect 15312 -14708 15408 -14692
rect 14319 -14760 15041 -14759
rect 14319 -15480 14320 -14760
rect 15040 -15480 15041 -14760
rect 14319 -15481 15041 -15480
rect 13900 -15548 13996 -15532
rect 15312 -15532 15328 -14708
rect 15392 -15532 15408 -14708
rect 16724 -14708 16820 -14692
rect 15731 -14760 16453 -14759
rect 15731 -15480 15732 -14760
rect 16452 -15480 16453 -14760
rect 15731 -15481 16453 -15480
rect 15312 -15548 15408 -15532
rect 16724 -15532 16740 -14708
rect 16804 -15532 16820 -14708
rect 18136 -14708 18232 -14692
rect 17143 -14760 17865 -14759
rect 17143 -15480 17144 -14760
rect 17864 -15480 17865 -14760
rect 17143 -15481 17865 -15480
rect 16724 -15548 16820 -15532
rect 18136 -15532 18152 -14708
rect 18216 -15532 18232 -14708
rect 19548 -14708 19644 -14692
rect 18555 -14760 19277 -14759
rect 18555 -15480 18556 -14760
rect 19276 -15480 19277 -14760
rect 18555 -15481 19277 -15480
rect 18136 -15548 18232 -15532
rect 19548 -15532 19564 -14708
rect 19628 -15532 19644 -14708
rect 20960 -14708 21056 -14692
rect 19967 -14760 20689 -14759
rect 19967 -15480 19968 -14760
rect 20688 -15480 20689 -14760
rect 19967 -15481 20689 -15480
rect 19548 -15548 19644 -15532
rect 20960 -15532 20976 -14708
rect 21040 -15532 21056 -14708
rect 22372 -14708 22468 -14692
rect 21379 -14760 22101 -14759
rect 21379 -15480 21380 -14760
rect 22100 -15480 22101 -14760
rect 21379 -15481 22101 -15480
rect 20960 -15548 21056 -15532
rect 22372 -15532 22388 -14708
rect 22452 -15532 22468 -14708
rect 23784 -14708 23880 -14692
rect 22791 -14760 23513 -14759
rect 22791 -15480 22792 -14760
rect 23512 -15480 23513 -14760
rect 22791 -15481 23513 -15480
rect 22372 -15548 22468 -15532
rect 23784 -15532 23800 -14708
rect 23864 -15532 23880 -14708
rect 23784 -15548 23880 -15532
rect -22812 -15828 -22716 -15812
rect -23805 -15880 -23083 -15879
rect -23805 -16600 -23804 -15880
rect -23084 -16600 -23083 -15880
rect -23805 -16601 -23083 -16600
rect -22812 -16652 -22796 -15828
rect -22732 -16652 -22716 -15828
rect -21400 -15828 -21304 -15812
rect -22393 -15880 -21671 -15879
rect -22393 -16600 -22392 -15880
rect -21672 -16600 -21671 -15880
rect -22393 -16601 -21671 -16600
rect -22812 -16668 -22716 -16652
rect -21400 -16652 -21384 -15828
rect -21320 -16652 -21304 -15828
rect -19988 -15828 -19892 -15812
rect -20981 -15880 -20259 -15879
rect -20981 -16600 -20980 -15880
rect -20260 -16600 -20259 -15880
rect -20981 -16601 -20259 -16600
rect -21400 -16668 -21304 -16652
rect -19988 -16652 -19972 -15828
rect -19908 -16652 -19892 -15828
rect -18576 -15828 -18480 -15812
rect -19569 -15880 -18847 -15879
rect -19569 -16600 -19568 -15880
rect -18848 -16600 -18847 -15880
rect -19569 -16601 -18847 -16600
rect -19988 -16668 -19892 -16652
rect -18576 -16652 -18560 -15828
rect -18496 -16652 -18480 -15828
rect -17164 -15828 -17068 -15812
rect -18157 -15880 -17435 -15879
rect -18157 -16600 -18156 -15880
rect -17436 -16600 -17435 -15880
rect -18157 -16601 -17435 -16600
rect -18576 -16668 -18480 -16652
rect -17164 -16652 -17148 -15828
rect -17084 -16652 -17068 -15828
rect -15752 -15828 -15656 -15812
rect -16745 -15880 -16023 -15879
rect -16745 -16600 -16744 -15880
rect -16024 -16600 -16023 -15880
rect -16745 -16601 -16023 -16600
rect -17164 -16668 -17068 -16652
rect -15752 -16652 -15736 -15828
rect -15672 -16652 -15656 -15828
rect -14340 -15828 -14244 -15812
rect -15333 -15880 -14611 -15879
rect -15333 -16600 -15332 -15880
rect -14612 -16600 -14611 -15880
rect -15333 -16601 -14611 -16600
rect -15752 -16668 -15656 -16652
rect -14340 -16652 -14324 -15828
rect -14260 -16652 -14244 -15828
rect -12928 -15828 -12832 -15812
rect -13921 -15880 -13199 -15879
rect -13921 -16600 -13920 -15880
rect -13200 -16600 -13199 -15880
rect -13921 -16601 -13199 -16600
rect -14340 -16668 -14244 -16652
rect -12928 -16652 -12912 -15828
rect -12848 -16652 -12832 -15828
rect -11516 -15828 -11420 -15812
rect -12509 -15880 -11787 -15879
rect -12509 -16600 -12508 -15880
rect -11788 -16600 -11787 -15880
rect -12509 -16601 -11787 -16600
rect -12928 -16668 -12832 -16652
rect -11516 -16652 -11500 -15828
rect -11436 -16652 -11420 -15828
rect -10104 -15828 -10008 -15812
rect -11097 -15880 -10375 -15879
rect -11097 -16600 -11096 -15880
rect -10376 -16600 -10375 -15880
rect -11097 -16601 -10375 -16600
rect -11516 -16668 -11420 -16652
rect -10104 -16652 -10088 -15828
rect -10024 -16652 -10008 -15828
rect -8692 -15828 -8596 -15812
rect -9685 -15880 -8963 -15879
rect -9685 -16600 -9684 -15880
rect -8964 -16600 -8963 -15880
rect -9685 -16601 -8963 -16600
rect -10104 -16668 -10008 -16652
rect -8692 -16652 -8676 -15828
rect -8612 -16652 -8596 -15828
rect -7280 -15828 -7184 -15812
rect -8273 -15880 -7551 -15879
rect -8273 -16600 -8272 -15880
rect -7552 -16600 -7551 -15880
rect -8273 -16601 -7551 -16600
rect -8692 -16668 -8596 -16652
rect -7280 -16652 -7264 -15828
rect -7200 -16652 -7184 -15828
rect -5868 -15828 -5772 -15812
rect -6861 -15880 -6139 -15879
rect -6861 -16600 -6860 -15880
rect -6140 -16600 -6139 -15880
rect -6861 -16601 -6139 -16600
rect -7280 -16668 -7184 -16652
rect -5868 -16652 -5852 -15828
rect -5788 -16652 -5772 -15828
rect -4456 -15828 -4360 -15812
rect -5449 -15880 -4727 -15879
rect -5449 -16600 -5448 -15880
rect -4728 -16600 -4727 -15880
rect -5449 -16601 -4727 -16600
rect -5868 -16668 -5772 -16652
rect -4456 -16652 -4440 -15828
rect -4376 -16652 -4360 -15828
rect -3044 -15828 -2948 -15812
rect -4037 -15880 -3315 -15879
rect -4037 -16600 -4036 -15880
rect -3316 -16600 -3315 -15880
rect -4037 -16601 -3315 -16600
rect -4456 -16668 -4360 -16652
rect -3044 -16652 -3028 -15828
rect -2964 -16652 -2948 -15828
rect -1632 -15828 -1536 -15812
rect -2625 -15880 -1903 -15879
rect -2625 -16600 -2624 -15880
rect -1904 -16600 -1903 -15880
rect -2625 -16601 -1903 -16600
rect -3044 -16668 -2948 -16652
rect -1632 -16652 -1616 -15828
rect -1552 -16652 -1536 -15828
rect -220 -15828 -124 -15812
rect -1213 -15880 -491 -15879
rect -1213 -16600 -1212 -15880
rect -492 -16600 -491 -15880
rect -1213 -16601 -491 -16600
rect -1632 -16668 -1536 -16652
rect -220 -16652 -204 -15828
rect -140 -16652 -124 -15828
rect 1192 -15828 1288 -15812
rect 199 -15880 921 -15879
rect 199 -16600 200 -15880
rect 920 -16600 921 -15880
rect 199 -16601 921 -16600
rect -220 -16668 -124 -16652
rect 1192 -16652 1208 -15828
rect 1272 -16652 1288 -15828
rect 2604 -15828 2700 -15812
rect 1611 -15880 2333 -15879
rect 1611 -16600 1612 -15880
rect 2332 -16600 2333 -15880
rect 1611 -16601 2333 -16600
rect 1192 -16668 1288 -16652
rect 2604 -16652 2620 -15828
rect 2684 -16652 2700 -15828
rect 4016 -15828 4112 -15812
rect 3023 -15880 3745 -15879
rect 3023 -16600 3024 -15880
rect 3744 -16600 3745 -15880
rect 3023 -16601 3745 -16600
rect 2604 -16668 2700 -16652
rect 4016 -16652 4032 -15828
rect 4096 -16652 4112 -15828
rect 5428 -15828 5524 -15812
rect 4435 -15880 5157 -15879
rect 4435 -16600 4436 -15880
rect 5156 -16600 5157 -15880
rect 4435 -16601 5157 -16600
rect 4016 -16668 4112 -16652
rect 5428 -16652 5444 -15828
rect 5508 -16652 5524 -15828
rect 6840 -15828 6936 -15812
rect 5847 -15880 6569 -15879
rect 5847 -16600 5848 -15880
rect 6568 -16600 6569 -15880
rect 5847 -16601 6569 -16600
rect 5428 -16668 5524 -16652
rect 6840 -16652 6856 -15828
rect 6920 -16652 6936 -15828
rect 8252 -15828 8348 -15812
rect 7259 -15880 7981 -15879
rect 7259 -16600 7260 -15880
rect 7980 -16600 7981 -15880
rect 7259 -16601 7981 -16600
rect 6840 -16668 6936 -16652
rect 8252 -16652 8268 -15828
rect 8332 -16652 8348 -15828
rect 9664 -15828 9760 -15812
rect 8671 -15880 9393 -15879
rect 8671 -16600 8672 -15880
rect 9392 -16600 9393 -15880
rect 8671 -16601 9393 -16600
rect 8252 -16668 8348 -16652
rect 9664 -16652 9680 -15828
rect 9744 -16652 9760 -15828
rect 11076 -15828 11172 -15812
rect 10083 -15880 10805 -15879
rect 10083 -16600 10084 -15880
rect 10804 -16600 10805 -15880
rect 10083 -16601 10805 -16600
rect 9664 -16668 9760 -16652
rect 11076 -16652 11092 -15828
rect 11156 -16652 11172 -15828
rect 12488 -15828 12584 -15812
rect 11495 -15880 12217 -15879
rect 11495 -16600 11496 -15880
rect 12216 -16600 12217 -15880
rect 11495 -16601 12217 -16600
rect 11076 -16668 11172 -16652
rect 12488 -16652 12504 -15828
rect 12568 -16652 12584 -15828
rect 13900 -15828 13996 -15812
rect 12907 -15880 13629 -15879
rect 12907 -16600 12908 -15880
rect 13628 -16600 13629 -15880
rect 12907 -16601 13629 -16600
rect 12488 -16668 12584 -16652
rect 13900 -16652 13916 -15828
rect 13980 -16652 13996 -15828
rect 15312 -15828 15408 -15812
rect 14319 -15880 15041 -15879
rect 14319 -16600 14320 -15880
rect 15040 -16600 15041 -15880
rect 14319 -16601 15041 -16600
rect 13900 -16668 13996 -16652
rect 15312 -16652 15328 -15828
rect 15392 -16652 15408 -15828
rect 16724 -15828 16820 -15812
rect 15731 -15880 16453 -15879
rect 15731 -16600 15732 -15880
rect 16452 -16600 16453 -15880
rect 15731 -16601 16453 -16600
rect 15312 -16668 15408 -16652
rect 16724 -16652 16740 -15828
rect 16804 -16652 16820 -15828
rect 18136 -15828 18232 -15812
rect 17143 -15880 17865 -15879
rect 17143 -16600 17144 -15880
rect 17864 -16600 17865 -15880
rect 17143 -16601 17865 -16600
rect 16724 -16668 16820 -16652
rect 18136 -16652 18152 -15828
rect 18216 -16652 18232 -15828
rect 19548 -15828 19644 -15812
rect 18555 -15880 19277 -15879
rect 18555 -16600 18556 -15880
rect 19276 -16600 19277 -15880
rect 18555 -16601 19277 -16600
rect 18136 -16668 18232 -16652
rect 19548 -16652 19564 -15828
rect 19628 -16652 19644 -15828
rect 20960 -15828 21056 -15812
rect 19967 -15880 20689 -15879
rect 19967 -16600 19968 -15880
rect 20688 -16600 20689 -15880
rect 19967 -16601 20689 -16600
rect 19548 -16668 19644 -16652
rect 20960 -16652 20976 -15828
rect 21040 -16652 21056 -15828
rect 22372 -15828 22468 -15812
rect 21379 -15880 22101 -15879
rect 21379 -16600 21380 -15880
rect 22100 -16600 22101 -15880
rect 21379 -16601 22101 -16600
rect 20960 -16668 21056 -16652
rect 22372 -16652 22388 -15828
rect 22452 -16652 22468 -15828
rect 23784 -15828 23880 -15812
rect 22791 -15880 23513 -15879
rect 22791 -16600 22792 -15880
rect 23512 -16600 23513 -15880
rect 22791 -16601 23513 -16600
rect 22372 -16668 22468 -16652
rect 23784 -16652 23800 -15828
rect 23864 -16652 23880 -15828
rect 23784 -16668 23880 -16652
rect -22812 -16948 -22716 -16932
rect -23805 -17000 -23083 -16999
rect -23805 -17720 -23804 -17000
rect -23084 -17720 -23083 -17000
rect -23805 -17721 -23083 -17720
rect -22812 -17772 -22796 -16948
rect -22732 -17772 -22716 -16948
rect -21400 -16948 -21304 -16932
rect -22393 -17000 -21671 -16999
rect -22393 -17720 -22392 -17000
rect -21672 -17720 -21671 -17000
rect -22393 -17721 -21671 -17720
rect -22812 -17788 -22716 -17772
rect -21400 -17772 -21384 -16948
rect -21320 -17772 -21304 -16948
rect -19988 -16948 -19892 -16932
rect -20981 -17000 -20259 -16999
rect -20981 -17720 -20980 -17000
rect -20260 -17720 -20259 -17000
rect -20981 -17721 -20259 -17720
rect -21400 -17788 -21304 -17772
rect -19988 -17772 -19972 -16948
rect -19908 -17772 -19892 -16948
rect -18576 -16948 -18480 -16932
rect -19569 -17000 -18847 -16999
rect -19569 -17720 -19568 -17000
rect -18848 -17720 -18847 -17000
rect -19569 -17721 -18847 -17720
rect -19988 -17788 -19892 -17772
rect -18576 -17772 -18560 -16948
rect -18496 -17772 -18480 -16948
rect -17164 -16948 -17068 -16932
rect -18157 -17000 -17435 -16999
rect -18157 -17720 -18156 -17000
rect -17436 -17720 -17435 -17000
rect -18157 -17721 -17435 -17720
rect -18576 -17788 -18480 -17772
rect -17164 -17772 -17148 -16948
rect -17084 -17772 -17068 -16948
rect -15752 -16948 -15656 -16932
rect -16745 -17000 -16023 -16999
rect -16745 -17720 -16744 -17000
rect -16024 -17720 -16023 -17000
rect -16745 -17721 -16023 -17720
rect -17164 -17788 -17068 -17772
rect -15752 -17772 -15736 -16948
rect -15672 -17772 -15656 -16948
rect -14340 -16948 -14244 -16932
rect -15333 -17000 -14611 -16999
rect -15333 -17720 -15332 -17000
rect -14612 -17720 -14611 -17000
rect -15333 -17721 -14611 -17720
rect -15752 -17788 -15656 -17772
rect -14340 -17772 -14324 -16948
rect -14260 -17772 -14244 -16948
rect -12928 -16948 -12832 -16932
rect -13921 -17000 -13199 -16999
rect -13921 -17720 -13920 -17000
rect -13200 -17720 -13199 -17000
rect -13921 -17721 -13199 -17720
rect -14340 -17788 -14244 -17772
rect -12928 -17772 -12912 -16948
rect -12848 -17772 -12832 -16948
rect -11516 -16948 -11420 -16932
rect -12509 -17000 -11787 -16999
rect -12509 -17720 -12508 -17000
rect -11788 -17720 -11787 -17000
rect -12509 -17721 -11787 -17720
rect -12928 -17788 -12832 -17772
rect -11516 -17772 -11500 -16948
rect -11436 -17772 -11420 -16948
rect -10104 -16948 -10008 -16932
rect -11097 -17000 -10375 -16999
rect -11097 -17720 -11096 -17000
rect -10376 -17720 -10375 -17000
rect -11097 -17721 -10375 -17720
rect -11516 -17788 -11420 -17772
rect -10104 -17772 -10088 -16948
rect -10024 -17772 -10008 -16948
rect -8692 -16948 -8596 -16932
rect -9685 -17000 -8963 -16999
rect -9685 -17720 -9684 -17000
rect -8964 -17720 -8963 -17000
rect -9685 -17721 -8963 -17720
rect -10104 -17788 -10008 -17772
rect -8692 -17772 -8676 -16948
rect -8612 -17772 -8596 -16948
rect -7280 -16948 -7184 -16932
rect -8273 -17000 -7551 -16999
rect -8273 -17720 -8272 -17000
rect -7552 -17720 -7551 -17000
rect -8273 -17721 -7551 -17720
rect -8692 -17788 -8596 -17772
rect -7280 -17772 -7264 -16948
rect -7200 -17772 -7184 -16948
rect -5868 -16948 -5772 -16932
rect -6861 -17000 -6139 -16999
rect -6861 -17720 -6860 -17000
rect -6140 -17720 -6139 -17000
rect -6861 -17721 -6139 -17720
rect -7280 -17788 -7184 -17772
rect -5868 -17772 -5852 -16948
rect -5788 -17772 -5772 -16948
rect -4456 -16948 -4360 -16932
rect -5449 -17000 -4727 -16999
rect -5449 -17720 -5448 -17000
rect -4728 -17720 -4727 -17000
rect -5449 -17721 -4727 -17720
rect -5868 -17788 -5772 -17772
rect -4456 -17772 -4440 -16948
rect -4376 -17772 -4360 -16948
rect -3044 -16948 -2948 -16932
rect -4037 -17000 -3315 -16999
rect -4037 -17720 -4036 -17000
rect -3316 -17720 -3315 -17000
rect -4037 -17721 -3315 -17720
rect -4456 -17788 -4360 -17772
rect -3044 -17772 -3028 -16948
rect -2964 -17772 -2948 -16948
rect -1632 -16948 -1536 -16932
rect -2625 -17000 -1903 -16999
rect -2625 -17720 -2624 -17000
rect -1904 -17720 -1903 -17000
rect -2625 -17721 -1903 -17720
rect -3044 -17788 -2948 -17772
rect -1632 -17772 -1616 -16948
rect -1552 -17772 -1536 -16948
rect -220 -16948 -124 -16932
rect -1213 -17000 -491 -16999
rect -1213 -17720 -1212 -17000
rect -492 -17720 -491 -17000
rect -1213 -17721 -491 -17720
rect -1632 -17788 -1536 -17772
rect -220 -17772 -204 -16948
rect -140 -17772 -124 -16948
rect 1192 -16948 1288 -16932
rect 199 -17000 921 -16999
rect 199 -17720 200 -17000
rect 920 -17720 921 -17000
rect 199 -17721 921 -17720
rect -220 -17788 -124 -17772
rect 1192 -17772 1208 -16948
rect 1272 -17772 1288 -16948
rect 2604 -16948 2700 -16932
rect 1611 -17000 2333 -16999
rect 1611 -17720 1612 -17000
rect 2332 -17720 2333 -17000
rect 1611 -17721 2333 -17720
rect 1192 -17788 1288 -17772
rect 2604 -17772 2620 -16948
rect 2684 -17772 2700 -16948
rect 4016 -16948 4112 -16932
rect 3023 -17000 3745 -16999
rect 3023 -17720 3024 -17000
rect 3744 -17720 3745 -17000
rect 3023 -17721 3745 -17720
rect 2604 -17788 2700 -17772
rect 4016 -17772 4032 -16948
rect 4096 -17772 4112 -16948
rect 5428 -16948 5524 -16932
rect 4435 -17000 5157 -16999
rect 4435 -17720 4436 -17000
rect 5156 -17720 5157 -17000
rect 4435 -17721 5157 -17720
rect 4016 -17788 4112 -17772
rect 5428 -17772 5444 -16948
rect 5508 -17772 5524 -16948
rect 6840 -16948 6936 -16932
rect 5847 -17000 6569 -16999
rect 5847 -17720 5848 -17000
rect 6568 -17720 6569 -17000
rect 5847 -17721 6569 -17720
rect 5428 -17788 5524 -17772
rect 6840 -17772 6856 -16948
rect 6920 -17772 6936 -16948
rect 8252 -16948 8348 -16932
rect 7259 -17000 7981 -16999
rect 7259 -17720 7260 -17000
rect 7980 -17720 7981 -17000
rect 7259 -17721 7981 -17720
rect 6840 -17788 6936 -17772
rect 8252 -17772 8268 -16948
rect 8332 -17772 8348 -16948
rect 9664 -16948 9760 -16932
rect 8671 -17000 9393 -16999
rect 8671 -17720 8672 -17000
rect 9392 -17720 9393 -17000
rect 8671 -17721 9393 -17720
rect 8252 -17788 8348 -17772
rect 9664 -17772 9680 -16948
rect 9744 -17772 9760 -16948
rect 11076 -16948 11172 -16932
rect 10083 -17000 10805 -16999
rect 10083 -17720 10084 -17000
rect 10804 -17720 10805 -17000
rect 10083 -17721 10805 -17720
rect 9664 -17788 9760 -17772
rect 11076 -17772 11092 -16948
rect 11156 -17772 11172 -16948
rect 12488 -16948 12584 -16932
rect 11495 -17000 12217 -16999
rect 11495 -17720 11496 -17000
rect 12216 -17720 12217 -17000
rect 11495 -17721 12217 -17720
rect 11076 -17788 11172 -17772
rect 12488 -17772 12504 -16948
rect 12568 -17772 12584 -16948
rect 13900 -16948 13996 -16932
rect 12907 -17000 13629 -16999
rect 12907 -17720 12908 -17000
rect 13628 -17720 13629 -17000
rect 12907 -17721 13629 -17720
rect 12488 -17788 12584 -17772
rect 13900 -17772 13916 -16948
rect 13980 -17772 13996 -16948
rect 15312 -16948 15408 -16932
rect 14319 -17000 15041 -16999
rect 14319 -17720 14320 -17000
rect 15040 -17720 15041 -17000
rect 14319 -17721 15041 -17720
rect 13900 -17788 13996 -17772
rect 15312 -17772 15328 -16948
rect 15392 -17772 15408 -16948
rect 16724 -16948 16820 -16932
rect 15731 -17000 16453 -16999
rect 15731 -17720 15732 -17000
rect 16452 -17720 16453 -17000
rect 15731 -17721 16453 -17720
rect 15312 -17788 15408 -17772
rect 16724 -17772 16740 -16948
rect 16804 -17772 16820 -16948
rect 18136 -16948 18232 -16932
rect 17143 -17000 17865 -16999
rect 17143 -17720 17144 -17000
rect 17864 -17720 17865 -17000
rect 17143 -17721 17865 -17720
rect 16724 -17788 16820 -17772
rect 18136 -17772 18152 -16948
rect 18216 -17772 18232 -16948
rect 19548 -16948 19644 -16932
rect 18555 -17000 19277 -16999
rect 18555 -17720 18556 -17000
rect 19276 -17720 19277 -17000
rect 18555 -17721 19277 -17720
rect 18136 -17788 18232 -17772
rect 19548 -17772 19564 -16948
rect 19628 -17772 19644 -16948
rect 20960 -16948 21056 -16932
rect 19967 -17000 20689 -16999
rect 19967 -17720 19968 -17000
rect 20688 -17720 20689 -17000
rect 19967 -17721 20689 -17720
rect 19548 -17788 19644 -17772
rect 20960 -17772 20976 -16948
rect 21040 -17772 21056 -16948
rect 22372 -16948 22468 -16932
rect 21379 -17000 22101 -16999
rect 21379 -17720 21380 -17000
rect 22100 -17720 22101 -17000
rect 21379 -17721 22101 -17720
rect 20960 -17788 21056 -17772
rect 22372 -17772 22388 -16948
rect 22452 -17772 22468 -16948
rect 23784 -16948 23880 -16932
rect 22791 -17000 23513 -16999
rect 22791 -17720 22792 -17000
rect 23512 -17720 23513 -17000
rect 22791 -17721 23513 -17720
rect 22372 -17788 22468 -17772
rect 23784 -17772 23800 -16948
rect 23864 -17772 23880 -16948
rect 23784 -17788 23880 -17772
rect -22812 -18068 -22716 -18052
rect -23805 -18120 -23083 -18119
rect -23805 -18840 -23804 -18120
rect -23084 -18840 -23083 -18120
rect -23805 -18841 -23083 -18840
rect -22812 -18892 -22796 -18068
rect -22732 -18892 -22716 -18068
rect -21400 -18068 -21304 -18052
rect -22393 -18120 -21671 -18119
rect -22393 -18840 -22392 -18120
rect -21672 -18840 -21671 -18120
rect -22393 -18841 -21671 -18840
rect -22812 -18908 -22716 -18892
rect -21400 -18892 -21384 -18068
rect -21320 -18892 -21304 -18068
rect -19988 -18068 -19892 -18052
rect -20981 -18120 -20259 -18119
rect -20981 -18840 -20980 -18120
rect -20260 -18840 -20259 -18120
rect -20981 -18841 -20259 -18840
rect -21400 -18908 -21304 -18892
rect -19988 -18892 -19972 -18068
rect -19908 -18892 -19892 -18068
rect -18576 -18068 -18480 -18052
rect -19569 -18120 -18847 -18119
rect -19569 -18840 -19568 -18120
rect -18848 -18840 -18847 -18120
rect -19569 -18841 -18847 -18840
rect -19988 -18908 -19892 -18892
rect -18576 -18892 -18560 -18068
rect -18496 -18892 -18480 -18068
rect -17164 -18068 -17068 -18052
rect -18157 -18120 -17435 -18119
rect -18157 -18840 -18156 -18120
rect -17436 -18840 -17435 -18120
rect -18157 -18841 -17435 -18840
rect -18576 -18908 -18480 -18892
rect -17164 -18892 -17148 -18068
rect -17084 -18892 -17068 -18068
rect -15752 -18068 -15656 -18052
rect -16745 -18120 -16023 -18119
rect -16745 -18840 -16744 -18120
rect -16024 -18840 -16023 -18120
rect -16745 -18841 -16023 -18840
rect -17164 -18908 -17068 -18892
rect -15752 -18892 -15736 -18068
rect -15672 -18892 -15656 -18068
rect -14340 -18068 -14244 -18052
rect -15333 -18120 -14611 -18119
rect -15333 -18840 -15332 -18120
rect -14612 -18840 -14611 -18120
rect -15333 -18841 -14611 -18840
rect -15752 -18908 -15656 -18892
rect -14340 -18892 -14324 -18068
rect -14260 -18892 -14244 -18068
rect -12928 -18068 -12832 -18052
rect -13921 -18120 -13199 -18119
rect -13921 -18840 -13920 -18120
rect -13200 -18840 -13199 -18120
rect -13921 -18841 -13199 -18840
rect -14340 -18908 -14244 -18892
rect -12928 -18892 -12912 -18068
rect -12848 -18892 -12832 -18068
rect -11516 -18068 -11420 -18052
rect -12509 -18120 -11787 -18119
rect -12509 -18840 -12508 -18120
rect -11788 -18840 -11787 -18120
rect -12509 -18841 -11787 -18840
rect -12928 -18908 -12832 -18892
rect -11516 -18892 -11500 -18068
rect -11436 -18892 -11420 -18068
rect -10104 -18068 -10008 -18052
rect -11097 -18120 -10375 -18119
rect -11097 -18840 -11096 -18120
rect -10376 -18840 -10375 -18120
rect -11097 -18841 -10375 -18840
rect -11516 -18908 -11420 -18892
rect -10104 -18892 -10088 -18068
rect -10024 -18892 -10008 -18068
rect -8692 -18068 -8596 -18052
rect -9685 -18120 -8963 -18119
rect -9685 -18840 -9684 -18120
rect -8964 -18840 -8963 -18120
rect -9685 -18841 -8963 -18840
rect -10104 -18908 -10008 -18892
rect -8692 -18892 -8676 -18068
rect -8612 -18892 -8596 -18068
rect -7280 -18068 -7184 -18052
rect -8273 -18120 -7551 -18119
rect -8273 -18840 -8272 -18120
rect -7552 -18840 -7551 -18120
rect -8273 -18841 -7551 -18840
rect -8692 -18908 -8596 -18892
rect -7280 -18892 -7264 -18068
rect -7200 -18892 -7184 -18068
rect -5868 -18068 -5772 -18052
rect -6861 -18120 -6139 -18119
rect -6861 -18840 -6860 -18120
rect -6140 -18840 -6139 -18120
rect -6861 -18841 -6139 -18840
rect -7280 -18908 -7184 -18892
rect -5868 -18892 -5852 -18068
rect -5788 -18892 -5772 -18068
rect -4456 -18068 -4360 -18052
rect -5449 -18120 -4727 -18119
rect -5449 -18840 -5448 -18120
rect -4728 -18840 -4727 -18120
rect -5449 -18841 -4727 -18840
rect -5868 -18908 -5772 -18892
rect -4456 -18892 -4440 -18068
rect -4376 -18892 -4360 -18068
rect -3044 -18068 -2948 -18052
rect -4037 -18120 -3315 -18119
rect -4037 -18840 -4036 -18120
rect -3316 -18840 -3315 -18120
rect -4037 -18841 -3315 -18840
rect -4456 -18908 -4360 -18892
rect -3044 -18892 -3028 -18068
rect -2964 -18892 -2948 -18068
rect -1632 -18068 -1536 -18052
rect -2625 -18120 -1903 -18119
rect -2625 -18840 -2624 -18120
rect -1904 -18840 -1903 -18120
rect -2625 -18841 -1903 -18840
rect -3044 -18908 -2948 -18892
rect -1632 -18892 -1616 -18068
rect -1552 -18892 -1536 -18068
rect -220 -18068 -124 -18052
rect -1213 -18120 -491 -18119
rect -1213 -18840 -1212 -18120
rect -492 -18840 -491 -18120
rect -1213 -18841 -491 -18840
rect -1632 -18908 -1536 -18892
rect -220 -18892 -204 -18068
rect -140 -18892 -124 -18068
rect 1192 -18068 1288 -18052
rect 199 -18120 921 -18119
rect 199 -18840 200 -18120
rect 920 -18840 921 -18120
rect 199 -18841 921 -18840
rect -220 -18908 -124 -18892
rect 1192 -18892 1208 -18068
rect 1272 -18892 1288 -18068
rect 2604 -18068 2700 -18052
rect 1611 -18120 2333 -18119
rect 1611 -18840 1612 -18120
rect 2332 -18840 2333 -18120
rect 1611 -18841 2333 -18840
rect 1192 -18908 1288 -18892
rect 2604 -18892 2620 -18068
rect 2684 -18892 2700 -18068
rect 4016 -18068 4112 -18052
rect 3023 -18120 3745 -18119
rect 3023 -18840 3024 -18120
rect 3744 -18840 3745 -18120
rect 3023 -18841 3745 -18840
rect 2604 -18908 2700 -18892
rect 4016 -18892 4032 -18068
rect 4096 -18892 4112 -18068
rect 5428 -18068 5524 -18052
rect 4435 -18120 5157 -18119
rect 4435 -18840 4436 -18120
rect 5156 -18840 5157 -18120
rect 4435 -18841 5157 -18840
rect 4016 -18908 4112 -18892
rect 5428 -18892 5444 -18068
rect 5508 -18892 5524 -18068
rect 6840 -18068 6936 -18052
rect 5847 -18120 6569 -18119
rect 5847 -18840 5848 -18120
rect 6568 -18840 6569 -18120
rect 5847 -18841 6569 -18840
rect 5428 -18908 5524 -18892
rect 6840 -18892 6856 -18068
rect 6920 -18892 6936 -18068
rect 8252 -18068 8348 -18052
rect 7259 -18120 7981 -18119
rect 7259 -18840 7260 -18120
rect 7980 -18840 7981 -18120
rect 7259 -18841 7981 -18840
rect 6840 -18908 6936 -18892
rect 8252 -18892 8268 -18068
rect 8332 -18892 8348 -18068
rect 9664 -18068 9760 -18052
rect 8671 -18120 9393 -18119
rect 8671 -18840 8672 -18120
rect 9392 -18840 9393 -18120
rect 8671 -18841 9393 -18840
rect 8252 -18908 8348 -18892
rect 9664 -18892 9680 -18068
rect 9744 -18892 9760 -18068
rect 11076 -18068 11172 -18052
rect 10083 -18120 10805 -18119
rect 10083 -18840 10084 -18120
rect 10804 -18840 10805 -18120
rect 10083 -18841 10805 -18840
rect 9664 -18908 9760 -18892
rect 11076 -18892 11092 -18068
rect 11156 -18892 11172 -18068
rect 12488 -18068 12584 -18052
rect 11495 -18120 12217 -18119
rect 11495 -18840 11496 -18120
rect 12216 -18840 12217 -18120
rect 11495 -18841 12217 -18840
rect 11076 -18908 11172 -18892
rect 12488 -18892 12504 -18068
rect 12568 -18892 12584 -18068
rect 13900 -18068 13996 -18052
rect 12907 -18120 13629 -18119
rect 12907 -18840 12908 -18120
rect 13628 -18840 13629 -18120
rect 12907 -18841 13629 -18840
rect 12488 -18908 12584 -18892
rect 13900 -18892 13916 -18068
rect 13980 -18892 13996 -18068
rect 15312 -18068 15408 -18052
rect 14319 -18120 15041 -18119
rect 14319 -18840 14320 -18120
rect 15040 -18840 15041 -18120
rect 14319 -18841 15041 -18840
rect 13900 -18908 13996 -18892
rect 15312 -18892 15328 -18068
rect 15392 -18892 15408 -18068
rect 16724 -18068 16820 -18052
rect 15731 -18120 16453 -18119
rect 15731 -18840 15732 -18120
rect 16452 -18840 16453 -18120
rect 15731 -18841 16453 -18840
rect 15312 -18908 15408 -18892
rect 16724 -18892 16740 -18068
rect 16804 -18892 16820 -18068
rect 18136 -18068 18232 -18052
rect 17143 -18120 17865 -18119
rect 17143 -18840 17144 -18120
rect 17864 -18840 17865 -18120
rect 17143 -18841 17865 -18840
rect 16724 -18908 16820 -18892
rect 18136 -18892 18152 -18068
rect 18216 -18892 18232 -18068
rect 19548 -18068 19644 -18052
rect 18555 -18120 19277 -18119
rect 18555 -18840 18556 -18120
rect 19276 -18840 19277 -18120
rect 18555 -18841 19277 -18840
rect 18136 -18908 18232 -18892
rect 19548 -18892 19564 -18068
rect 19628 -18892 19644 -18068
rect 20960 -18068 21056 -18052
rect 19967 -18120 20689 -18119
rect 19967 -18840 19968 -18120
rect 20688 -18840 20689 -18120
rect 19967 -18841 20689 -18840
rect 19548 -18908 19644 -18892
rect 20960 -18892 20976 -18068
rect 21040 -18892 21056 -18068
rect 22372 -18068 22468 -18052
rect 21379 -18120 22101 -18119
rect 21379 -18840 21380 -18120
rect 22100 -18840 22101 -18120
rect 21379 -18841 22101 -18840
rect 20960 -18908 21056 -18892
rect 22372 -18892 22388 -18068
rect 22452 -18892 22468 -18068
rect 23784 -18068 23880 -18052
rect 22791 -18120 23513 -18119
rect 22791 -18840 22792 -18120
rect 23512 -18840 23513 -18120
rect 22791 -18841 23513 -18840
rect 22372 -18908 22468 -18892
rect 23784 -18892 23800 -18068
rect 23864 -18892 23880 -18068
rect 23784 -18908 23880 -18892
<< properties >>
string FIXED_BBOX 22712 18040 23592 18920
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4 l 4 val 35.04 carea 2.00 cperi 0.19 nx 34 ny 34 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
