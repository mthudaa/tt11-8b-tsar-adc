magic
tech sky130A
magscale 1 2
timestamp 1746260845
<< nwell >>
rect -246 -4435 246 4435
<< pmos >>
rect -50 3916 50 4216
rect -50 3488 50 3788
rect -50 3060 50 3360
rect -50 2632 50 2932
rect -50 2204 50 2504
rect -50 1776 50 2076
rect -50 1348 50 1648
rect -50 920 50 1220
rect -50 492 50 792
rect -50 64 50 364
rect -50 -364 50 -64
rect -50 -792 50 -492
rect -50 -1220 50 -920
rect -50 -1648 50 -1348
rect -50 -2076 50 -1776
rect -50 -2504 50 -2204
rect -50 -2932 50 -2632
rect -50 -3360 50 -3060
rect -50 -3788 50 -3488
rect -50 -4216 50 -3916
<< pdiff >>
rect -108 4204 -50 4216
rect -108 3928 -96 4204
rect -62 3928 -50 4204
rect -108 3916 -50 3928
rect 50 4204 108 4216
rect 50 3928 62 4204
rect 96 3928 108 4204
rect 50 3916 108 3928
rect -108 3776 -50 3788
rect -108 3500 -96 3776
rect -62 3500 -50 3776
rect -108 3488 -50 3500
rect 50 3776 108 3788
rect 50 3500 62 3776
rect 96 3500 108 3776
rect 50 3488 108 3500
rect -108 3348 -50 3360
rect -108 3072 -96 3348
rect -62 3072 -50 3348
rect -108 3060 -50 3072
rect 50 3348 108 3360
rect 50 3072 62 3348
rect 96 3072 108 3348
rect 50 3060 108 3072
rect -108 2920 -50 2932
rect -108 2644 -96 2920
rect -62 2644 -50 2920
rect -108 2632 -50 2644
rect 50 2920 108 2932
rect 50 2644 62 2920
rect 96 2644 108 2920
rect 50 2632 108 2644
rect -108 2492 -50 2504
rect -108 2216 -96 2492
rect -62 2216 -50 2492
rect -108 2204 -50 2216
rect 50 2492 108 2504
rect 50 2216 62 2492
rect 96 2216 108 2492
rect 50 2204 108 2216
rect -108 2064 -50 2076
rect -108 1788 -96 2064
rect -62 1788 -50 2064
rect -108 1776 -50 1788
rect 50 2064 108 2076
rect 50 1788 62 2064
rect 96 1788 108 2064
rect 50 1776 108 1788
rect -108 1636 -50 1648
rect -108 1360 -96 1636
rect -62 1360 -50 1636
rect -108 1348 -50 1360
rect 50 1636 108 1648
rect 50 1360 62 1636
rect 96 1360 108 1636
rect 50 1348 108 1360
rect -108 1208 -50 1220
rect -108 932 -96 1208
rect -62 932 -50 1208
rect -108 920 -50 932
rect 50 1208 108 1220
rect 50 932 62 1208
rect 96 932 108 1208
rect 50 920 108 932
rect -108 780 -50 792
rect -108 504 -96 780
rect -62 504 -50 780
rect -108 492 -50 504
rect 50 780 108 792
rect 50 504 62 780
rect 96 504 108 780
rect 50 492 108 504
rect -108 352 -50 364
rect -108 76 -96 352
rect -62 76 -50 352
rect -108 64 -50 76
rect 50 352 108 364
rect 50 76 62 352
rect 96 76 108 352
rect 50 64 108 76
rect -108 -76 -50 -64
rect -108 -352 -96 -76
rect -62 -352 -50 -76
rect -108 -364 -50 -352
rect 50 -76 108 -64
rect 50 -352 62 -76
rect 96 -352 108 -76
rect 50 -364 108 -352
rect -108 -504 -50 -492
rect -108 -780 -96 -504
rect -62 -780 -50 -504
rect -108 -792 -50 -780
rect 50 -504 108 -492
rect 50 -780 62 -504
rect 96 -780 108 -504
rect 50 -792 108 -780
rect -108 -932 -50 -920
rect -108 -1208 -96 -932
rect -62 -1208 -50 -932
rect -108 -1220 -50 -1208
rect 50 -932 108 -920
rect 50 -1208 62 -932
rect 96 -1208 108 -932
rect 50 -1220 108 -1208
rect -108 -1360 -50 -1348
rect -108 -1636 -96 -1360
rect -62 -1636 -50 -1360
rect -108 -1648 -50 -1636
rect 50 -1360 108 -1348
rect 50 -1636 62 -1360
rect 96 -1636 108 -1360
rect 50 -1648 108 -1636
rect -108 -1788 -50 -1776
rect -108 -2064 -96 -1788
rect -62 -2064 -50 -1788
rect -108 -2076 -50 -2064
rect 50 -1788 108 -1776
rect 50 -2064 62 -1788
rect 96 -2064 108 -1788
rect 50 -2076 108 -2064
rect -108 -2216 -50 -2204
rect -108 -2492 -96 -2216
rect -62 -2492 -50 -2216
rect -108 -2504 -50 -2492
rect 50 -2216 108 -2204
rect 50 -2492 62 -2216
rect 96 -2492 108 -2216
rect 50 -2504 108 -2492
rect -108 -2644 -50 -2632
rect -108 -2920 -96 -2644
rect -62 -2920 -50 -2644
rect -108 -2932 -50 -2920
rect 50 -2644 108 -2632
rect 50 -2920 62 -2644
rect 96 -2920 108 -2644
rect 50 -2932 108 -2920
rect -108 -3072 -50 -3060
rect -108 -3348 -96 -3072
rect -62 -3348 -50 -3072
rect -108 -3360 -50 -3348
rect 50 -3072 108 -3060
rect 50 -3348 62 -3072
rect 96 -3348 108 -3072
rect 50 -3360 108 -3348
rect -108 -3500 -50 -3488
rect -108 -3776 -96 -3500
rect -62 -3776 -50 -3500
rect -108 -3788 -50 -3776
rect 50 -3500 108 -3488
rect 50 -3776 62 -3500
rect 96 -3776 108 -3500
rect 50 -3788 108 -3776
rect -108 -3928 -50 -3916
rect -108 -4204 -96 -3928
rect -62 -4204 -50 -3928
rect -108 -4216 -50 -4204
rect 50 -3928 108 -3916
rect 50 -4204 62 -3928
rect 96 -4204 108 -3928
rect 50 -4216 108 -4204
<< pdiffc >>
rect -96 3928 -62 4204
rect 62 3928 96 4204
rect -96 3500 -62 3776
rect 62 3500 96 3776
rect -96 3072 -62 3348
rect 62 3072 96 3348
rect -96 2644 -62 2920
rect 62 2644 96 2920
rect -96 2216 -62 2492
rect 62 2216 96 2492
rect -96 1788 -62 2064
rect 62 1788 96 2064
rect -96 1360 -62 1636
rect 62 1360 96 1636
rect -96 932 -62 1208
rect 62 932 96 1208
rect -96 504 -62 780
rect 62 504 96 780
rect -96 76 -62 352
rect 62 76 96 352
rect -96 -352 -62 -76
rect 62 -352 96 -76
rect -96 -780 -62 -504
rect 62 -780 96 -504
rect -96 -1208 -62 -932
rect 62 -1208 96 -932
rect -96 -1636 -62 -1360
rect 62 -1636 96 -1360
rect -96 -2064 -62 -1788
rect 62 -2064 96 -1788
rect -96 -2492 -62 -2216
rect 62 -2492 96 -2216
rect -96 -2920 -62 -2644
rect 62 -2920 96 -2644
rect -96 -3348 -62 -3072
rect 62 -3348 96 -3072
rect -96 -3776 -62 -3500
rect 62 -3776 96 -3500
rect -96 -4204 -62 -3928
rect 62 -4204 96 -3928
<< nsubdiff >>
rect -210 4365 -114 4399
rect 114 4365 210 4399
rect -210 4303 -176 4365
rect 176 4303 210 4365
rect -210 -4365 -176 -4303
rect 176 -4365 210 -4303
rect -210 -4399 -114 -4365
rect 114 -4399 210 -4365
<< nsubdiffcont >>
rect -114 4365 114 4399
rect -210 -4303 -176 4303
rect 176 -4303 210 4303
rect -114 -4399 114 -4365
<< poly >>
rect -50 4297 50 4313
rect -50 4263 -34 4297
rect 34 4263 50 4297
rect -50 4216 50 4263
rect -50 3869 50 3916
rect -50 3835 -34 3869
rect 34 3835 50 3869
rect -50 3788 50 3835
rect -50 3441 50 3488
rect -50 3407 -34 3441
rect 34 3407 50 3441
rect -50 3360 50 3407
rect -50 3013 50 3060
rect -50 2979 -34 3013
rect 34 2979 50 3013
rect -50 2932 50 2979
rect -50 2585 50 2632
rect -50 2551 -34 2585
rect 34 2551 50 2585
rect -50 2504 50 2551
rect -50 2157 50 2204
rect -50 2123 -34 2157
rect 34 2123 50 2157
rect -50 2076 50 2123
rect -50 1729 50 1776
rect -50 1695 -34 1729
rect 34 1695 50 1729
rect -50 1648 50 1695
rect -50 1301 50 1348
rect -50 1267 -34 1301
rect 34 1267 50 1301
rect -50 1220 50 1267
rect -50 873 50 920
rect -50 839 -34 873
rect 34 839 50 873
rect -50 792 50 839
rect -50 445 50 492
rect -50 411 -34 445
rect 34 411 50 445
rect -50 364 50 411
rect -50 17 50 64
rect -50 -17 -34 17
rect 34 -17 50 17
rect -50 -64 50 -17
rect -50 -411 50 -364
rect -50 -445 -34 -411
rect 34 -445 50 -411
rect -50 -492 50 -445
rect -50 -839 50 -792
rect -50 -873 -34 -839
rect 34 -873 50 -839
rect -50 -920 50 -873
rect -50 -1267 50 -1220
rect -50 -1301 -34 -1267
rect 34 -1301 50 -1267
rect -50 -1348 50 -1301
rect -50 -1695 50 -1648
rect -50 -1729 -34 -1695
rect 34 -1729 50 -1695
rect -50 -1776 50 -1729
rect -50 -2123 50 -2076
rect -50 -2157 -34 -2123
rect 34 -2157 50 -2123
rect -50 -2204 50 -2157
rect -50 -2551 50 -2504
rect -50 -2585 -34 -2551
rect 34 -2585 50 -2551
rect -50 -2632 50 -2585
rect -50 -2979 50 -2932
rect -50 -3013 -34 -2979
rect 34 -3013 50 -2979
rect -50 -3060 50 -3013
rect -50 -3407 50 -3360
rect -50 -3441 -34 -3407
rect 34 -3441 50 -3407
rect -50 -3488 50 -3441
rect -50 -3835 50 -3788
rect -50 -3869 -34 -3835
rect 34 -3869 50 -3835
rect -50 -3916 50 -3869
rect -50 -4263 50 -4216
rect -50 -4297 -34 -4263
rect 34 -4297 50 -4263
rect -50 -4313 50 -4297
<< polycont >>
rect -34 4263 34 4297
rect -34 3835 34 3869
rect -34 3407 34 3441
rect -34 2979 34 3013
rect -34 2551 34 2585
rect -34 2123 34 2157
rect -34 1695 34 1729
rect -34 1267 34 1301
rect -34 839 34 873
rect -34 411 34 445
rect -34 -17 34 17
rect -34 -445 34 -411
rect -34 -873 34 -839
rect -34 -1301 34 -1267
rect -34 -1729 34 -1695
rect -34 -2157 34 -2123
rect -34 -2585 34 -2551
rect -34 -3013 34 -2979
rect -34 -3441 34 -3407
rect -34 -3869 34 -3835
rect -34 -4297 34 -4263
<< locali >>
rect -210 4365 -114 4399
rect 114 4365 210 4399
rect -210 4303 -176 4365
rect 176 4303 210 4365
rect -50 4263 -34 4297
rect 34 4263 50 4297
rect -96 4204 -62 4220
rect -96 3912 -62 3928
rect 62 4204 96 4220
rect 62 3912 96 3928
rect -50 3835 -34 3869
rect 34 3835 50 3869
rect -96 3776 -62 3792
rect -96 3484 -62 3500
rect 62 3776 96 3792
rect 62 3484 96 3500
rect -50 3407 -34 3441
rect 34 3407 50 3441
rect -96 3348 -62 3364
rect -96 3056 -62 3072
rect 62 3348 96 3364
rect 62 3056 96 3072
rect -50 2979 -34 3013
rect 34 2979 50 3013
rect -96 2920 -62 2936
rect -96 2628 -62 2644
rect 62 2920 96 2936
rect 62 2628 96 2644
rect -50 2551 -34 2585
rect 34 2551 50 2585
rect -96 2492 -62 2508
rect -96 2200 -62 2216
rect 62 2492 96 2508
rect 62 2200 96 2216
rect -50 2123 -34 2157
rect 34 2123 50 2157
rect -96 2064 -62 2080
rect -96 1772 -62 1788
rect 62 2064 96 2080
rect 62 1772 96 1788
rect -50 1695 -34 1729
rect 34 1695 50 1729
rect -96 1636 -62 1652
rect -96 1344 -62 1360
rect 62 1636 96 1652
rect 62 1344 96 1360
rect -50 1267 -34 1301
rect 34 1267 50 1301
rect -96 1208 -62 1224
rect -96 916 -62 932
rect 62 1208 96 1224
rect 62 916 96 932
rect -50 839 -34 873
rect 34 839 50 873
rect -96 780 -62 796
rect -96 488 -62 504
rect 62 780 96 796
rect 62 488 96 504
rect -50 411 -34 445
rect 34 411 50 445
rect -96 352 -62 368
rect -96 60 -62 76
rect 62 352 96 368
rect 62 60 96 76
rect -50 -17 -34 17
rect 34 -17 50 17
rect -96 -76 -62 -60
rect -96 -368 -62 -352
rect 62 -76 96 -60
rect 62 -368 96 -352
rect -50 -445 -34 -411
rect 34 -445 50 -411
rect -96 -504 -62 -488
rect -96 -796 -62 -780
rect 62 -504 96 -488
rect 62 -796 96 -780
rect -50 -873 -34 -839
rect 34 -873 50 -839
rect -96 -932 -62 -916
rect -96 -1224 -62 -1208
rect 62 -932 96 -916
rect 62 -1224 96 -1208
rect -50 -1301 -34 -1267
rect 34 -1301 50 -1267
rect -96 -1360 -62 -1344
rect -96 -1652 -62 -1636
rect 62 -1360 96 -1344
rect 62 -1652 96 -1636
rect -50 -1729 -34 -1695
rect 34 -1729 50 -1695
rect -96 -1788 -62 -1772
rect -96 -2080 -62 -2064
rect 62 -1788 96 -1772
rect 62 -2080 96 -2064
rect -50 -2157 -34 -2123
rect 34 -2157 50 -2123
rect -96 -2216 -62 -2200
rect -96 -2508 -62 -2492
rect 62 -2216 96 -2200
rect 62 -2508 96 -2492
rect -50 -2585 -34 -2551
rect 34 -2585 50 -2551
rect -96 -2644 -62 -2628
rect -96 -2936 -62 -2920
rect 62 -2644 96 -2628
rect 62 -2936 96 -2920
rect -50 -3013 -34 -2979
rect 34 -3013 50 -2979
rect -96 -3072 -62 -3056
rect -96 -3364 -62 -3348
rect 62 -3072 96 -3056
rect 62 -3364 96 -3348
rect -50 -3441 -34 -3407
rect 34 -3441 50 -3407
rect -96 -3500 -62 -3484
rect -96 -3792 -62 -3776
rect 62 -3500 96 -3484
rect 62 -3792 96 -3776
rect -50 -3869 -34 -3835
rect 34 -3869 50 -3835
rect -96 -3928 -62 -3912
rect -96 -4220 -62 -4204
rect 62 -3928 96 -3912
rect 62 -4220 96 -4204
rect -50 -4297 -34 -4263
rect 34 -4297 50 -4263
rect -210 -4365 -176 -4303
rect 176 -4365 210 -4303
rect -210 -4399 -114 -4365
rect 114 -4399 210 -4365
<< viali >>
rect -34 4263 34 4297
rect -96 3928 -62 4204
rect 62 3928 96 4204
rect -34 3835 34 3869
rect -96 3500 -62 3776
rect 62 3500 96 3776
rect -34 3407 34 3441
rect -96 3072 -62 3348
rect 62 3072 96 3348
rect -34 2979 34 3013
rect -96 2644 -62 2920
rect 62 2644 96 2920
rect -34 2551 34 2585
rect -96 2216 -62 2492
rect 62 2216 96 2492
rect -34 2123 34 2157
rect -96 1788 -62 2064
rect 62 1788 96 2064
rect -34 1695 34 1729
rect -96 1360 -62 1636
rect 62 1360 96 1636
rect -34 1267 34 1301
rect -96 932 -62 1208
rect 62 932 96 1208
rect -34 839 34 873
rect -96 504 -62 780
rect 62 504 96 780
rect -34 411 34 445
rect -96 76 -62 352
rect 62 76 96 352
rect -34 -17 34 17
rect -96 -352 -62 -76
rect 62 -352 96 -76
rect -34 -445 34 -411
rect -96 -780 -62 -504
rect 62 -780 96 -504
rect -34 -873 34 -839
rect -96 -1208 -62 -932
rect 62 -1208 96 -932
rect -34 -1301 34 -1267
rect -96 -1636 -62 -1360
rect 62 -1636 96 -1360
rect -34 -1729 34 -1695
rect -96 -2064 -62 -1788
rect 62 -2064 96 -1788
rect -34 -2157 34 -2123
rect -96 -2492 -62 -2216
rect 62 -2492 96 -2216
rect -34 -2585 34 -2551
rect -96 -2920 -62 -2644
rect 62 -2920 96 -2644
rect -34 -3013 34 -2979
rect -96 -3348 -62 -3072
rect 62 -3348 96 -3072
rect -34 -3441 34 -3407
rect -96 -3776 -62 -3500
rect 62 -3776 96 -3500
rect -34 -3869 34 -3835
rect -96 -4204 -62 -3928
rect 62 -4204 96 -3928
rect -34 -4297 34 -4263
<< metal1 >>
rect -46 4297 46 4303
rect -46 4263 -34 4297
rect 34 4263 46 4297
rect -46 4257 46 4263
rect -102 4204 -56 4216
rect -102 3928 -96 4204
rect -62 3928 -56 4204
rect -102 3916 -56 3928
rect 56 4204 102 4216
rect 56 3928 62 4204
rect 96 3928 102 4204
rect 56 3916 102 3928
rect -46 3869 46 3875
rect -46 3835 -34 3869
rect 34 3835 46 3869
rect -46 3829 46 3835
rect -102 3776 -56 3788
rect -102 3500 -96 3776
rect -62 3500 -56 3776
rect -102 3488 -56 3500
rect 56 3776 102 3788
rect 56 3500 62 3776
rect 96 3500 102 3776
rect 56 3488 102 3500
rect -46 3441 46 3447
rect -46 3407 -34 3441
rect 34 3407 46 3441
rect -46 3401 46 3407
rect -102 3348 -56 3360
rect -102 3072 -96 3348
rect -62 3072 -56 3348
rect -102 3060 -56 3072
rect 56 3348 102 3360
rect 56 3072 62 3348
rect 96 3072 102 3348
rect 56 3060 102 3072
rect -46 3013 46 3019
rect -46 2979 -34 3013
rect 34 2979 46 3013
rect -46 2973 46 2979
rect -102 2920 -56 2932
rect -102 2644 -96 2920
rect -62 2644 -56 2920
rect -102 2632 -56 2644
rect 56 2920 102 2932
rect 56 2644 62 2920
rect 96 2644 102 2920
rect 56 2632 102 2644
rect -46 2585 46 2591
rect -46 2551 -34 2585
rect 34 2551 46 2585
rect -46 2545 46 2551
rect -102 2492 -56 2504
rect -102 2216 -96 2492
rect -62 2216 -56 2492
rect -102 2204 -56 2216
rect 56 2492 102 2504
rect 56 2216 62 2492
rect 96 2216 102 2492
rect 56 2204 102 2216
rect -46 2157 46 2163
rect -46 2123 -34 2157
rect 34 2123 46 2157
rect -46 2117 46 2123
rect -102 2064 -56 2076
rect -102 1788 -96 2064
rect -62 1788 -56 2064
rect -102 1776 -56 1788
rect 56 2064 102 2076
rect 56 1788 62 2064
rect 96 1788 102 2064
rect 56 1776 102 1788
rect -46 1729 46 1735
rect -46 1695 -34 1729
rect 34 1695 46 1729
rect -46 1689 46 1695
rect -102 1636 -56 1648
rect -102 1360 -96 1636
rect -62 1360 -56 1636
rect -102 1348 -56 1360
rect 56 1636 102 1648
rect 56 1360 62 1636
rect 96 1360 102 1636
rect 56 1348 102 1360
rect -46 1301 46 1307
rect -46 1267 -34 1301
rect 34 1267 46 1301
rect -46 1261 46 1267
rect -102 1208 -56 1220
rect -102 932 -96 1208
rect -62 932 -56 1208
rect -102 920 -56 932
rect 56 1208 102 1220
rect 56 932 62 1208
rect 96 932 102 1208
rect 56 920 102 932
rect -46 873 46 879
rect -46 839 -34 873
rect 34 839 46 873
rect -46 833 46 839
rect -102 780 -56 792
rect -102 504 -96 780
rect -62 504 -56 780
rect -102 492 -56 504
rect 56 780 102 792
rect 56 504 62 780
rect 96 504 102 780
rect 56 492 102 504
rect -46 445 46 451
rect -46 411 -34 445
rect 34 411 46 445
rect -46 405 46 411
rect -102 352 -56 364
rect -102 76 -96 352
rect -62 76 -56 352
rect -102 64 -56 76
rect 56 352 102 364
rect 56 76 62 352
rect 96 76 102 352
rect 56 64 102 76
rect -46 17 46 23
rect -46 -17 -34 17
rect 34 -17 46 17
rect -46 -23 46 -17
rect -102 -76 -56 -64
rect -102 -352 -96 -76
rect -62 -352 -56 -76
rect -102 -364 -56 -352
rect 56 -76 102 -64
rect 56 -352 62 -76
rect 96 -352 102 -76
rect 56 -364 102 -352
rect -46 -411 46 -405
rect -46 -445 -34 -411
rect 34 -445 46 -411
rect -46 -451 46 -445
rect -102 -504 -56 -492
rect -102 -780 -96 -504
rect -62 -780 -56 -504
rect -102 -792 -56 -780
rect 56 -504 102 -492
rect 56 -780 62 -504
rect 96 -780 102 -504
rect 56 -792 102 -780
rect -46 -839 46 -833
rect -46 -873 -34 -839
rect 34 -873 46 -839
rect -46 -879 46 -873
rect -102 -932 -56 -920
rect -102 -1208 -96 -932
rect -62 -1208 -56 -932
rect -102 -1220 -56 -1208
rect 56 -932 102 -920
rect 56 -1208 62 -932
rect 96 -1208 102 -932
rect 56 -1220 102 -1208
rect -46 -1267 46 -1261
rect -46 -1301 -34 -1267
rect 34 -1301 46 -1267
rect -46 -1307 46 -1301
rect -102 -1360 -56 -1348
rect -102 -1636 -96 -1360
rect -62 -1636 -56 -1360
rect -102 -1648 -56 -1636
rect 56 -1360 102 -1348
rect 56 -1636 62 -1360
rect 96 -1636 102 -1360
rect 56 -1648 102 -1636
rect -46 -1695 46 -1689
rect -46 -1729 -34 -1695
rect 34 -1729 46 -1695
rect -46 -1735 46 -1729
rect -102 -1788 -56 -1776
rect -102 -2064 -96 -1788
rect -62 -2064 -56 -1788
rect -102 -2076 -56 -2064
rect 56 -1788 102 -1776
rect 56 -2064 62 -1788
rect 96 -2064 102 -1788
rect 56 -2076 102 -2064
rect -46 -2123 46 -2117
rect -46 -2157 -34 -2123
rect 34 -2157 46 -2123
rect -46 -2163 46 -2157
rect -102 -2216 -56 -2204
rect -102 -2492 -96 -2216
rect -62 -2492 -56 -2216
rect -102 -2504 -56 -2492
rect 56 -2216 102 -2204
rect 56 -2492 62 -2216
rect 96 -2492 102 -2216
rect 56 -2504 102 -2492
rect -46 -2551 46 -2545
rect -46 -2585 -34 -2551
rect 34 -2585 46 -2551
rect -46 -2591 46 -2585
rect -102 -2644 -56 -2632
rect -102 -2920 -96 -2644
rect -62 -2920 -56 -2644
rect -102 -2932 -56 -2920
rect 56 -2644 102 -2632
rect 56 -2920 62 -2644
rect 96 -2920 102 -2644
rect 56 -2932 102 -2920
rect -46 -2979 46 -2973
rect -46 -3013 -34 -2979
rect 34 -3013 46 -2979
rect -46 -3019 46 -3013
rect -102 -3072 -56 -3060
rect -102 -3348 -96 -3072
rect -62 -3348 -56 -3072
rect -102 -3360 -56 -3348
rect 56 -3072 102 -3060
rect 56 -3348 62 -3072
rect 96 -3348 102 -3072
rect 56 -3360 102 -3348
rect -46 -3407 46 -3401
rect -46 -3441 -34 -3407
rect 34 -3441 46 -3407
rect -46 -3447 46 -3441
rect -102 -3500 -56 -3488
rect -102 -3776 -96 -3500
rect -62 -3776 -56 -3500
rect -102 -3788 -56 -3776
rect 56 -3500 102 -3488
rect 56 -3776 62 -3500
rect 96 -3776 102 -3500
rect 56 -3788 102 -3776
rect -46 -3835 46 -3829
rect -46 -3869 -34 -3835
rect 34 -3869 46 -3835
rect -46 -3875 46 -3869
rect -102 -3928 -56 -3916
rect -102 -4204 -96 -3928
rect -62 -4204 -56 -3928
rect -102 -4216 -56 -4204
rect 56 -3928 102 -3916
rect 56 -4204 62 -3928
rect 96 -4204 102 -3928
rect 56 -4216 102 -4204
rect -46 -4263 46 -4257
rect -46 -4297 -34 -4263
rect 34 -4297 46 -4263
rect -46 -4303 46 -4297
<< properties >>
string FIXED_BBOX -193 -4382 193 4382
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.5 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
