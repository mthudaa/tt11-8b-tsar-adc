magic
tech sky130A
magscale 1 2
timestamp 1746183267
<< viali >>
rect -17 369 6213 403
rect 6285 -17 9463 17
<< metal1 >>
rect -53 403 9499 439
rect -53 369 -17 403
rect 6213 369 9499 403
rect -53 363 9499 369
rect -53 289 9289 323
rect -53 143 119 243
rect 9327 143 9499 243
rect 166 63 9499 97
rect -53 17 9499 23
rect -53 -17 6285 17
rect 9463 -17 9499 17
rect -53 -53 9499 -17
use sky130_fd_pr__pfet_01v8_D9Q956  XM1
timestamp 1746182548
transform 0 1 3098 -1 0 193
box -246 -3151 246 3151
use sky130_fd_pr__nfet_01v8_H9ZN2D  XM2
timestamp 1746182548
transform 0 1 7874 -1 0 193
box -246 -1625 246 1625
<< labels >>
flabel metal1 -32 391 -15 407 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 -33 -34 -16 -18 0 FreeSans 400 0 0 0 VSS
port 1 nsew
flabel metal1 -43 300 -26 316 0 FreeSans 400 0 0 0 IN
port 2 nsew
flabel metal1 -42 184 -25 200 0 FreeSans 400 0 0 0 SWP
port 3 nsew
flabel metal1 9472 178 9490 195 0 FreeSans 400 0 0 0 SWN
port 4 nsew
flabel metal1 9474 73 9492 90 0 FreeSans 400 0 0 0 OUT
port 6 nsew
<< end >>
