magic
tech sky130A
magscale 1 2
timestamp 1747692869
<< metal1 >>
rect -22832 -34710 -22822 -34606
rect -22718 -34710 -18586 -34606
rect -18482 -34710 -18472 -34606
rect -25656 -34923 -25646 -34819
rect -25542 -34923 -17174 -34819
rect -17070 -34923 -17060 -34819
rect -28480 -35131 -28470 -35027
rect -28366 -35131 -14350 -35027
rect -14246 -35131 -14236 -35027
rect -34128 -35338 -34118 -35234
rect -34014 -35338 -8702 -35234
rect -8598 -35338 -8588 -35234
rect -45174 -36038 -20206 -35934
rect -20102 -36038 2594 -35934
rect -45174 -36246 -21170 -36142
rect -21066 -36246 2594 -36142
rect -45174 -36454 -22478 -36350
rect -22374 -36454 2594 -36350
rect -45174 -36662 -21618 -36558
rect -21514 -36662 2594 -36558
rect -45174 -36870 -22686 -36766
rect -22582 -36870 2594 -36766
rect -45174 -37078 -19998 -36974
rect -19894 -37078 2594 -36974
rect -45174 -37286 -21410 -37182
rect -21306 -37286 2594 -37182
rect -45174 -37494 -18586 -37390
rect -18482 -37494 2594 -37390
rect -45174 -37702 -17174 -37598
rect -17070 -37702 2594 -37598
rect -45174 -37910 -28470 -37806
rect -28366 -37910 2594 -37806
rect -45174 -38118 -8702 -38014
rect -8598 -38118 2594 -38014
<< via1 >>
rect -22822 -34710 -22718 -34606
rect -18586 -34710 -18482 -34606
rect -25646 -34923 -25542 -34819
rect -17174 -34923 -17070 -34819
rect -28470 -35131 -28366 -35027
rect -14350 -35131 -14246 -35027
rect -34118 -35338 -34014 -35234
rect -8702 -35338 -8598 -35234
rect -20206 -36038 -20102 -35934
rect -21170 -36246 -21066 -36142
rect -22478 -36454 -22374 -36350
rect -21618 -36662 -21514 -36558
rect -22686 -36870 -22582 -36766
rect -19998 -37078 -19894 -36974
rect -21410 -37286 -21306 -37182
rect -18586 -37494 -18482 -37390
rect -17174 -37702 -17070 -37598
rect -28470 -37910 -28366 -37806
rect -8702 -38118 -8598 -38014
<< metal2 >>
rect -21410 -7726 -21306 -7716
rect -22686 -14446 -22582 -14436
rect -22686 -21166 -22582 -14550
rect -21618 -15566 -21514 -15556
rect -34118 -34606 -34014 -34596
rect -34118 -35234 -34014 -34710
rect -34118 -35349 -34014 -35338
rect -28470 -34606 -28366 -34596
rect -28470 -35027 -28366 -34710
rect -25646 -34606 -25542 -34596
rect -25646 -34819 -25542 -34710
rect -22822 -34606 -22718 -34596
rect -22822 -34720 -22718 -34710
rect -25646 -34933 -25542 -34923
rect -28470 -37806 -28366 -35131
rect -22686 -36766 -22582 -21270
rect -22478 -16926 -22374 -16916
rect -22478 -36350 -22374 -17030
rect -22478 -36464 -22374 -36454
rect -21618 -18926 -21514 -15670
rect -21618 -36558 -21514 -19030
rect -21618 -36672 -21514 -36662
rect -21410 -34606 -21306 -7830
rect -19998 -12206 -19894 -12196
rect -20206 -16686 -20102 -16676
rect -22686 -36880 -22582 -36870
rect -21410 -37182 -21306 -34710
rect -21170 -16926 -21066 -16916
rect -21170 -36142 -21066 -17030
rect -20206 -35934 -20102 -16790
rect -20206 -36048 -20102 -36038
rect -19998 -25646 -19894 -12310
rect -21170 -36256 -21066 -36246
rect -19998 -36974 -19894 -25750
rect -19998 -37088 -19894 -37078
rect -18586 -34606 -18482 -34596
rect -21410 -37296 -21306 -37286
rect -18586 -37390 -18482 -34710
rect -18586 -37504 -18482 -37494
rect -17174 -34606 -17070 -34596
rect -17174 -34819 -17070 -34710
rect -17174 -37598 -17070 -34923
rect -14350 -34606 -14246 -34596
rect -14350 -35027 -14246 -34710
rect -14350 -35141 -14246 -35131
rect -8702 -34606 -8598 -34596
rect -17174 -37712 -17070 -37702
rect -8702 -35234 -8598 -34710
rect -28470 -37920 -28366 -37910
rect -8702 -38014 -8598 -35338
rect -8702 -38128 -8598 -38118
<< via2 >>
rect -21410 -7830 -21306 -7726
rect -22686 -14550 -22582 -14446
rect -21618 -15670 -21514 -15566
rect -22686 -21270 -22582 -21166
rect -34118 -34710 -34014 -34606
rect -28470 -34710 -28366 -34606
rect -25646 -34710 -25542 -34606
rect -22822 -34710 -22718 -34606
rect -22478 -17030 -22374 -16926
rect -21618 -19030 -21514 -18926
rect -19998 -12310 -19894 -12206
rect -20206 -16790 -20102 -16686
rect -21410 -34710 -21306 -34606
rect -21170 -17030 -21066 -16926
rect -19998 -25750 -19894 -25646
rect -18586 -34710 -18482 -34606
rect -17174 -34710 -17070 -34606
rect -14350 -34710 -14246 -34606
rect -8702 -34710 -8598 -34606
<< metal3 >>
rect -43762 -34606 -32706 891
rect -43762 -34710 -34118 -34606
rect -34014 -34710 -32706 -34606
rect -32466 -34606 -27058 890
rect -32466 -34710 -28470 -34606
rect -28366 -34710 -27058 -34606
rect -26818 -34606 -24233 890
rect -26818 -34710 -25646 -34606
rect -25542 -34710 -24233 -34606
rect -23994 -34601 -22822 890
rect -22583 -7726 -19997 891
rect -22583 -7830 -21410 -7726
rect -21306 -7830 -19997 -7726
rect -22583 -7831 -19997 -7830
rect -21420 -7835 -21296 -7831
rect -22582 -12201 -19998 -8070
rect -22582 -12206 -19884 -12201
rect -22582 -12310 -19998 -12206
rect -19894 -12310 -19884 -12206
rect -20008 -12315 -19884 -12310
rect -22582 -14441 -19998 -12550
rect -22696 -14446 -19998 -14441
rect -22696 -14550 -22686 -14446
rect -22582 -14550 -19998 -14446
rect -22696 -14555 -19998 -14550
rect -22582 -15566 -19998 -14790
rect -22582 -15670 -21618 -15566
rect -21514 -15670 -19998 -15566
rect -21628 -15675 -21504 -15670
rect -22582 -16926 -21410 -15910
rect -20216 -16686 -20092 -16681
rect -20216 -16790 -20206 -16686
rect -20102 -16790 -20092 -16686
rect -20216 -16795 -20092 -16790
rect -22582 -17030 -22478 -16926
rect -22374 -17030 -21410 -16926
rect -22582 -17910 -21410 -17030
rect -21180 -16926 -21056 -16921
rect -21180 -17030 -21170 -16926
rect -21066 -17030 -21056 -16926
rect -21180 -17035 -21056 -17030
rect -22582 -18926 -19998 -18150
rect -22582 -19030 -21618 -18926
rect -21514 -19030 -19998 -18926
rect -21628 -19035 -21504 -19030
rect -22582 -21161 -19999 -19270
rect -22696 -21166 -19999 -21161
rect -22696 -21270 -22686 -21166
rect -22582 -21270 -19999 -21166
rect -22696 -21275 -19999 -21270
rect -22582 -25641 -19998 -21510
rect -22582 -25646 -19884 -25641
rect -22582 -25750 -19998 -25646
rect -19894 -25750 -19884 -25646
rect -20008 -25755 -19884 -25750
rect -23994 -34606 -22708 -34601
rect -23994 -34710 -22822 -34606
rect -22718 -34710 -22708 -34606
rect -22582 -34606 -19996 -25988
rect -22582 -34710 -21410 -34606
rect -21306 -34710 -19996 -34606
rect -19758 -34601 -18586 890
rect -19758 -34606 -18472 -34601
rect -19758 -34710 -18586 -34606
rect -18482 -34710 -18472 -34606
rect -18347 -34606 -15762 890
rect -18347 -34710 -17174 -34606
rect -17070 -34710 -15762 -34606
rect -15522 -34606 -10114 890
rect -15522 -34710 -14350 -34606
rect -14246 -34710 -10114 -34606
rect -9874 -34606 1182 890
rect -9874 -34710 -8702 -34606
rect -8598 -34710 1182 -34606
rect -34128 -34715 -34004 -34710
rect -28480 -34715 -28356 -34710
rect -25656 -34715 -25532 -34710
rect -22832 -34715 -22708 -34710
rect -21420 -34715 -21296 -34710
rect -18596 -34715 -18472 -34710
rect -17184 -34715 -17060 -34710
rect -14360 -34715 -14236 -34710
rect -9874 -34711 1182 -34710
rect -8712 -34715 -8588 -34711
<< metal4 >>
rect -43683 1209 811 1931
rect -43683 -34631 -42961 1209
rect -42271 -34631 -41549 1209
rect -40859 -34631 -40137 1209
rect -39447 -34631 -38725 1209
rect -38035 -34631 -37313 1209
rect -36623 -34631 -35901 1209
rect -35211 -34631 -34489 1209
rect -33799 -34631 -33077 1209
rect -32387 -34631 -31665 1209
rect -30975 -34631 -30253 1209
rect -29563 -34631 -28841 1209
rect -28151 -34631 -27429 1209
rect -26739 -34631 -26017 1209
rect -25327 -34631 -24605 1209
rect -23915 -34631 -23193 1209
rect -22503 -34631 -21781 1209
rect -21091 -34631 -20369 1209
rect -19679 -34631 -18957 1209
rect -18267 -34631 -17545 1209
rect -16855 -34631 -16133 1209
rect -15443 -34631 -14721 1209
rect -14031 -34631 -13309 1209
rect -12619 -34631 -11897 1209
rect -11207 -34631 -10485 1209
rect -9795 -34631 -9073 1209
rect -8383 -34631 -7661 1209
rect -6971 -34631 -6249 1209
rect -5559 -34631 -4837 1209
rect -4147 -34631 -3425 1209
rect -2735 -34631 -2013 1209
rect -1323 -34631 -601 1209
rect 89 -34631 811 1209
use sky130_fd_pr__cap_mim_m3_1_8CZEMF  sky130_fd_pr__cap_mim_m3_1_8CZEMF_0
timestamp 1747692682
transform 1 0 -21290 0 1 -17470
box -23884 -18360 23884 18360
<< labels >>
flabel metal1 -45174 -36038 -20206 -35934 0 FreeSans 800 0 0 0 VCM
port 0 nsew
flabel metal1 -45174 -36246 -21170 -36142 0 FreeSans 800 0 0 0 SW[9]
port 1 nsew
flabel metal1 -45174 -36454 -22478 -36350 0 FreeSans 800 0 0 0 SW[8]
port 2 nsew
flabel metal1 -45174 -36662 -21618 -36558 0 FreeSans 800 0 0 0 SW[7]
port 3 nsew
flabel metal1 -45174 -36870 -22686 -36766 0 FreeSans 800 0 0 0 SW[6]
port 4 nsew
flabel metal1 -45174 -37078 -19998 -36974 0 FreeSans 800 0 0 0 SW[5]
port 5 nsew
flabel metal1 -45174 -37286 -21410 -37182 0 FreeSans 800 0 0 0 SW[4]
port 6 nsew
flabel metal1 -45174 -37494 -18586 -37390 0 FreeSans 800 0 0 0 SW[3]
port 7 nsew
flabel metal1 -45174 -37702 -17174 -37598 0 FreeSans 800 0 0 0 SW[2]
port 8 nsew
flabel metal1 -45174 -37910 -28470 -37806 0 FreeSans 800 0 0 0 SW[1]
port 9 nsew
flabel metal1 -45174 -38118 -8702 -38014 0 FreeSans 800 0 0 0 SW[0]
port 10 nsew
flabel metal4 -43683 1209 811 1931 0 FreeSans 800 0 0 0 VC
port 14 nsew
<< end >>
