magic
tech sky130A
magscale 1 2
timestamp 1746262095
<< viali >>
rect 142 1527 8940 1561
rect 142 -123 4580 -89
<< metal1 >>
rect 106 1561 8976 1597
rect 106 1527 142 1561
rect 8940 1527 8976 1561
rect 106 1521 8976 1527
rect 325 1447 8757 1521
rect 106 1301 176 1401
rect 228 1301 284 1401
rect 337 1061 8757 1255
rect 106 915 284 1015
rect 106 569 8976 869
rect 106 423 284 523
rect 316 183 4406 377
rect 166 37 176 137
rect 228 37 284 137
rect 316 -83 4406 -9
rect 106 -89 8976 -83
rect 106 -123 142 -89
rect 4580 -123 8976 -89
rect 106 -159 8976 -123
<< via1 >>
rect 176 1301 228 1401
rect 176 37 228 137
<< metal2 >>
rect 176 1401 228 1411
rect 176 137 228 1301
rect 176 27 228 37
use sky130_fd_pr__nfet_01v8_MKNP2D  sky130_fd_pr__nfet_01v8_MKNP2D_0
timestamp 1746260845
transform 0 1 2361 -1 0 87
box -246 -2255 246 2255
use sky130_fd_pr__pfet_01v8_C9QZQZ  sky130_fd_pr__pfet_01v8_C9QZQZ_0
timestamp 1746260845
transform 0 1 4541 -1 0 965
box -246 -4435 246 4435
use sky130_fd_pr__pfet_01v8_C9QZQZ  XM1
timestamp 1746260845
transform 0 1 4541 -1 0 1351
box -246 -4435 246 4435
use sky130_fd_pr__nfet_01v8_MKNP2D  XM3
timestamp 1746260845
transform 0 1 2361 -1 0 473
box -246 -2255 246 2255
<< labels >>
flabel metal1 120 1555 128 1563 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 117 1345 122 1350 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 120 961 125 966 0 FreeSans 400 0 0 0 CKB
port 2 nsew
flabel metal1 120 469 125 474 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel metal1 122 -124 127 -119 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 8943 715 8948 720 0 FreeSans 400 0 0 0 OUT
port 6 nsew
<< end >>
