magic
tech sky130A
magscale 1 2
timestamp 1747656850
<< viali >>
rect 238 1527 1996 1561
rect 238 -123 1124 -89
<< metal1 >>
rect 106 1561 2128 1597
rect 106 1527 238 1561
rect 1996 1527 2128 1561
rect 106 1521 2128 1527
rect 325 1447 1909 1521
rect 106 1301 176 1401
rect 228 1301 283 1401
rect 325 1061 1909 1255
rect 106 915 284 1015
rect 106 570 2128 869
rect 106 423 284 523
rect 316 183 1046 377
rect 166 37 176 137
rect 228 37 284 137
rect 316 -83 1046 -9
rect 106 -89 2128 -83
rect 106 -123 238 -89
rect 1124 -123 2128 -89
rect 106 -159 2128 -123
<< via1 >>
rect 176 1301 228 1401
rect 176 37 228 137
<< metal2 >>
rect 176 1401 228 1411
rect 176 137 228 1301
rect 176 27 228 37
use sky130_fd_pr__nfet_01v8_KT5VMN  sky130_fd_pr__nfet_01v8_KT5VMN_0
timestamp 1747652019
transform 0 1 681 -1 0 87
box -246 -575 246 575
use sky130_fd_pr__pfet_01v8_NMYCWJ  sky130_fd_pr__pfet_01v8_NMYCWJ_0
timestamp 1747652019
transform 0 1 1117 -1 0 965
box -246 -1011 246 1011
use sky130_fd_pr__pfet_01v8_NMYCWJ  XM1
timestamp 1747652019
transform 0 1 1117 -1 0 1351
box -246 -1011 246 1011
use sky130_fd_pr__nfet_01v8_KT5VMN  XM3
timestamp 1747652019
transform 0 1 681 -1 0 473
box -246 -575 246 575
<< labels >>
flabel metal1 106 1521 238 1597 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 106 1301 176 1401 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 106 915 284 1015 0 FreeSans 400 0 0 0 CKB
port 2 nsew
flabel metal1 106 423 284 523 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel metal1 106 -159 238 -83 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 1962 666 2074 747 0 FreeSans 400 0 0 0 OUT
port 6 nsew
<< end >>
