magic
tech sky130A
magscale 1 2
timestamp 1747524117
<< viali >>
rect 238 1527 3708 1561
rect 238 -123 1964 -89
<< metal1 >>
rect 106 1561 3840 1597
rect 106 1527 238 1561
rect 3708 1527 3840 1561
rect 106 1521 3840 1527
rect 325 1447 3621 1521
rect 106 1301 176 1401
rect 228 1301 284 1401
rect 325 1061 3621 1255
rect 106 915 284 1015
rect 106 569 3840 868
rect 106 423 284 523
rect 316 183 1886 377
rect 166 37 176 137
rect 228 37 280 137
rect 316 -83 1886 -9
rect 106 -89 3840 -83
rect 106 -123 238 -89
rect 1964 -123 3840 -89
rect 106 -159 3840 -123
<< via1 >>
rect 176 1301 228 1401
rect 176 37 228 137
<< metal2 >>
rect 176 1401 228 1411
rect 176 137 228 1301
rect 176 27 228 37
use sky130_fd_pr__nfet_01v8_X73VMN  sky130_fd_pr__nfet_01v8_X73VMN_0
timestamp 1747524117
transform 0 1 1101 -1 0 87
box -246 -995 246 995
use sky130_fd_pr__pfet_01v8_NMYLRJ  sky130_fd_pr__pfet_01v8_NMYLRJ_0
timestamp 1747524117
transform 0 1 1973 -1 0 965
box -246 -1867 246 1867
use sky130_fd_pr__pfet_01v8_NMYLRJ  XM1
timestamp 1747524117
transform 0 1 1973 -1 0 1351
box -246 -1867 246 1867
use sky130_fd_pr__nfet_01v8_X73VMN  XM3
timestamp 1747524117
transform 0 1 1101 -1 0 473
box -246 -995 246 995
<< labels >>
flabel metal1 106 1521 238 1597 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 106 1301 176 1401 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 106 915 284 1015 0 FreeSans 400 0 0 0 CKB
port 2 nsew
flabel metal1 106 423 284 523 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel metal1 106 -159 238 -83 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 3667 678 3799 754 0 FreeSans 400 0 0 0 OUT
port 6 nsew
<< end >>
