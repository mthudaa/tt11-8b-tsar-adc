magic
tech sky130A
magscale 1 2
timestamp 1746259868
<< pwell >>
rect -246 -575 246 575
<< nmos >>
rect -50 265 50 365
rect -50 55 50 155
rect -50 -155 50 -55
rect -50 -365 50 -265
<< ndiff >>
rect -108 353 -50 365
rect -108 277 -96 353
rect -62 277 -50 353
rect -108 265 -50 277
rect 50 353 108 365
rect 50 277 62 353
rect 96 277 108 353
rect 50 265 108 277
rect -108 143 -50 155
rect -108 67 -96 143
rect -62 67 -50 143
rect -108 55 -50 67
rect 50 143 108 155
rect 50 67 62 143
rect 96 67 108 143
rect 50 55 108 67
rect -108 -67 -50 -55
rect -108 -143 -96 -67
rect -62 -143 -50 -67
rect -108 -155 -50 -143
rect 50 -67 108 -55
rect 50 -143 62 -67
rect 96 -143 108 -67
rect 50 -155 108 -143
rect -108 -277 -50 -265
rect -108 -353 -96 -277
rect -62 -353 -50 -277
rect -108 -365 -50 -353
rect 50 -277 108 -265
rect 50 -353 62 -277
rect 96 -353 108 -277
rect 50 -365 108 -353
<< ndiffc >>
rect -96 277 -62 353
rect 62 277 96 353
rect -96 67 -62 143
rect 62 67 96 143
rect -96 -143 -62 -67
rect 62 -143 96 -67
rect -96 -353 -62 -277
rect 62 -353 96 -277
<< psubdiff >>
rect -210 505 -114 539
rect 114 505 210 539
rect -210 443 -176 505
rect 176 443 210 505
rect -210 -505 -176 -443
rect 176 -505 210 -443
rect -210 -539 -114 -505
rect 114 -539 210 -505
<< psubdiffcont >>
rect -114 505 114 539
rect -210 -443 -176 443
rect 176 -443 210 443
rect -114 -539 114 -505
<< poly >>
rect -50 437 50 453
rect -50 403 -34 437
rect 34 403 50 437
rect -50 365 50 403
rect -50 227 50 265
rect -50 193 -34 227
rect 34 193 50 227
rect -50 155 50 193
rect -50 17 50 55
rect -50 -17 -34 17
rect 34 -17 50 17
rect -50 -55 50 -17
rect -50 -193 50 -155
rect -50 -227 -34 -193
rect 34 -227 50 -193
rect -50 -265 50 -227
rect -50 -403 50 -365
rect -50 -437 -34 -403
rect 34 -437 50 -403
rect -50 -453 50 -437
<< polycont >>
rect -34 403 34 437
rect -34 193 34 227
rect -34 -17 34 17
rect -34 -227 34 -193
rect -34 -437 34 -403
<< locali >>
rect -210 505 -114 539
rect 114 505 210 539
rect -210 443 -176 505
rect 176 443 210 505
rect -50 403 -34 437
rect 34 403 50 437
rect -96 353 -62 369
rect -96 261 -62 277
rect 62 353 96 369
rect 62 261 96 277
rect -50 193 -34 227
rect 34 193 50 227
rect -96 143 -62 159
rect -96 51 -62 67
rect 62 143 96 159
rect 62 51 96 67
rect -50 -17 -34 17
rect 34 -17 50 17
rect -96 -67 -62 -51
rect -96 -159 -62 -143
rect 62 -67 96 -51
rect 62 -159 96 -143
rect -50 -227 -34 -193
rect 34 -227 50 -193
rect -96 -277 -62 -261
rect -96 -369 -62 -353
rect 62 -277 96 -261
rect 62 -369 96 -353
rect -50 -437 -34 -403
rect 34 -437 50 -403
rect -210 -505 -176 -443
rect 176 -505 210 -443
rect -210 -539 -114 -505
rect 114 -539 210 -505
<< viali >>
rect -34 403 34 437
rect -96 277 -62 353
rect 62 277 96 353
rect -34 193 34 227
rect -96 67 -62 143
rect 62 67 96 143
rect -34 -17 34 17
rect -96 -143 -62 -67
rect 62 -143 96 -67
rect -34 -227 34 -193
rect -96 -353 -62 -277
rect 62 -353 96 -277
rect -34 -437 34 -403
<< metal1 >>
rect -46 437 46 443
rect -46 403 -34 437
rect 34 403 46 437
rect -46 397 46 403
rect -102 353 -56 365
rect -102 277 -96 353
rect -62 277 -56 353
rect -102 265 -56 277
rect 56 353 102 365
rect 56 277 62 353
rect 96 277 102 353
rect 56 265 102 277
rect -46 227 46 233
rect -46 193 -34 227
rect 34 193 46 227
rect -46 187 46 193
rect -102 143 -56 155
rect -102 67 -96 143
rect -62 67 -56 143
rect -102 55 -56 67
rect 56 143 102 155
rect 56 67 62 143
rect 96 67 102 143
rect 56 55 102 67
rect -46 17 46 23
rect -46 -17 -34 17
rect 34 -17 46 17
rect -46 -23 46 -17
rect -102 -67 -56 -55
rect -102 -143 -96 -67
rect -62 -143 -56 -67
rect -102 -155 -56 -143
rect 56 -67 102 -55
rect 56 -143 62 -67
rect 96 -143 102 -67
rect 56 -155 102 -143
rect -46 -193 46 -187
rect -46 -227 -34 -193
rect 34 -227 46 -193
rect -46 -233 46 -227
rect -102 -277 -56 -265
rect -102 -353 -96 -277
rect -62 -353 -56 -277
rect -102 -365 -56 -353
rect 56 -277 102 -265
rect 56 -353 62 -277
rect 96 -353 102 -277
rect 56 -365 102 -353
rect -46 -403 46 -397
rect -46 -437 -34 -403
rect 34 -437 46 -403
rect -46 -443 46 -437
<< properties >>
string FIXED_BBOX -193 -522 193 522
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.5 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
