* NGSPICE file created from sar8b.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_2 abstract view
.subckt sky130_fd_sc_hs__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hs__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfrtp_1 abstract view
.subckt sky130_fd_sc_hs__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_8 abstract view
.subckt sky130_fd_sc_hs__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_1 abstract view
.subckt sky130_fd_sc_hs__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfxtp_1 abstract view
.subckt sky130_fd_sc_hs__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__decap_4 abstract view
.subckt sky130_fd_sc_hs__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_1 abstract view
.subckt sky130_fd_sc_hs__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfrtp_2 abstract view
.subckt sky130_fd_sc_hs__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor2_1 abstract view
.subckt sky130_fd_sc_hs__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and2_1 abstract view
.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_16 abstract view
.subckt sky130_fd_sc_hs__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__a21bo_1 abstract view
.subckt sky130_fd_sc_hs__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__o21a_1 abstract view
.subckt sky130_fd_sc_hs__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__or3b_1 abstract view
.subckt sky130_fd_sc_hs__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nand2_1 abstract view
.subckt sky130_fd_sc_hs__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__or4bb_1 abstract view
.subckt sky130_fd_sc_hs__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_2 abstract view
.subckt sky130_fd_sc_hs__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__buf_1 abstract view
.subckt sky130_fd_sc_hs__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_8 abstract view
.subckt sky130_fd_sc_hs__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__buf_2 abstract view
.subckt sky130_fd_sc_hs__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfxtp_4 abstract view
.subckt sky130_fd_sc_hs__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__o211a_1 abstract view
.subckt sky130_fd_sc_hs__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and3_1 abstract view
.subckt sky130_fd_sc_hs__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__xor2_1 abstract view
.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor3_1 abstract view
.subckt sky130_fd_sc_hs__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

.subckt sar8b CF[0] CF[1] CF[2] CF[3] CF[4] CF[5] CF[6] CF[7] CKO CKS CKSB CLK CMP_N
+ CMP_P DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] EN RDY SWN[0]
+ SWN[1] SWN[2] SWN[3] SWN[4] SWN[5] SWN[6] SWN[7] SWP[0] SWP[1] SWP[2] SWP[3] SWP[4]
+ SWP[5] SWP[6] SWP[7] VGND VPWR
XFILLER_0_11_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_8_55 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_66_ net6 net1 net14 VGND VGND VPWR VPWR net25 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_49_ clknet_1_0__leaf_CLK _03_ VGND VGND VPWR VPWR clk_div_0.COUNT\[1\] sky130_fd_sc_hs__dfxtp_1
XFILLER_0_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput31 net31 VGND VGND VPWR VPWR SWN[7] sky130_fd_sc_hs__clkbuf_1
Xoutput20 net20 VGND VGND VPWR VPWR DATA[4] sky130_fd_sc_hs__clkbuf_1
Xoutput7 net7 VGND VGND VPWR VPWR CF[2] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_65_ net7 net1 net14 VGND VGND VPWR VPWR net26 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_48_ clknet_1_0__leaf_CLK _02_ VGND VGND VPWR VPWR clk_div_0.COUNT\[0\] sky130_fd_sc_hs__dfxtp_1
XPHY_EDGE_ROW_8_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
Xoutput21 net21 VGND VGND VPWR VPWR DATA[5] sky130_fd_sc_hs__clkbuf_1
Xoutput32 net32 VGND VGND VPWR VPWR SWP[0] sky130_fd_sc_hs__clkbuf_1
Xoutput8 net8 VGND VGND VPWR VPWR CF[3] sky130_fd_sc_hs__clkbuf_1
Xoutput10 net10 VGND VGND VPWR VPWR CF[5] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_64_ net8 net1 net14 VGND VGND VPWR VPWR net27 sky130_fd_sc_hs__dfrtp_1
X_47_ net4 net12 net14 VGND VGND VPWR VPWR cyclic_flag_0.FINAL sky130_fd_sc_hs__dfrtp_2
XFILLER_0_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
Xoutput22 net22 VGND VGND VPWR VPWR DATA[6] sky130_fd_sc_hs__clkbuf_1
Xoutput33 net33 VGND VGND VPWR VPWR SWP[1] sky130_fd_sc_hs__clkbuf_1
Xoutput9 net9 VGND VGND VPWR VPWR CF[4] sky130_fd_sc_hs__clkbuf_1
Xoutput11 net11 VGND VGND VPWR VPWR CF[6] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_63_ net9 net1 net14 VGND VGND VPWR VPWR net28 sky130_fd_sc_hs__dfrtp_1
X_46_ net4 net11 net14 VGND VGND VPWR VPWR net12 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_5_48 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_29_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] VGND VGND VPWR VPWR _13_ sky130_fd_sc_hs__nor2_1
XFILLER_0_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_15_68 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput23 net23 VGND VGND VPWR VPWR DATA[7] sky130_fd_sc_hs__clkbuf_1
Xoutput12 net12 VGND VGND VPWR VPWR CF[7] sky130_fd_sc_hs__clkbuf_1
Xoutput34 net34 VGND VGND VPWR VPWR SWP[2] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_62_ net10 net1 net14 VGND VGND VPWR VPWR net29 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_45_ net4 net10 net14 VGND VGND VPWR VPWR net11 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_5_49 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_28_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] VGND VGND VPWR VPWR _12_ sky130_fd_sc_hs__and2_1
XTAP_TAPCELL_ROW_15_69 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
Xoutput24 net24 VGND VGND VPWR VPWR SWN[0] sky130_fd_sc_hs__clkbuf_1
Xoutput13 net13 VGND VGND VPWR VPWR CKO sky130_fd_sc_hs__clkbuf_1
Xoutput35 net35 VGND VGND VPWR VPWR SWP[3] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_61_ net11 net1 net14 VGND VGND VPWR VPWR net30 sky130_fd_sc_hs__dfrtp_1
Xclkbuf_1_1__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_1__leaf_CLK sky130_fd_sc_hs__clkbuf_16
XFILLER_0_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_44_ net4 net9 net14 VGND VGND VPWR VPWR net10 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_27_ clk_div_0.COUNT\[0\] _08_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hs__nor2_1
Xoutput25 net25 VGND VGND VPWR VPWR SWN[1] sky130_fd_sc_hs__clkbuf_1
Xoutput14 net14 VGND VGND VPWR VPWR CKS sky130_fd_sc_hs__clkbuf_1
Xoutput36 net36 VGND VGND VPWR VPWR SWP[4] sky130_fd_sc_hs__clkbuf_1
XPHY_EDGE_ROW_15_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_0_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_60_ net12 net1 net14 VGND VGND VPWR VPWR net31 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_43_ net4 net8 net14 VGND VGND VPWR VPWR net9 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_3_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_26_ _11_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_6_50 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xoutput26 net26 VGND VGND VPWR VPWR SWN[2] sky130_fd_sc_hs__clkbuf_1
Xoutput37 net37 VGND VGND VPWR VPWR SWP[5] sky130_fd_sc_hs__clkbuf_1
Xoutput15 net15 VGND VGND VPWR VPWR CKSB sky130_fd_sc_hs__clkbuf_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_16_70 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_7_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_42_ net4 net7 net14 VGND VGND VPWR VPWR net8 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_25_ net14 _10_ _09_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hs__a21bo_1
XTAP_TAPCELL_ROW_6_51 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
Xoutput16 net16 VGND VGND VPWR VPWR DATA[0] sky130_fd_sc_hs__clkbuf_1
Xoutput27 net27 VGND VGND VPWR VPWR SWN[3] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_9_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
Xoutput38 net38 VGND VGND VPWR VPWR SWP[6] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_16_71 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_41_ net4 net6 net14 VGND VGND VPWR VPWR net7 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_24_ net3 _07_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hs__and2_1
XFILLER_0_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
Xoutput17 net17 VGND VGND VPWR VPWR DATA[1] sky130_fd_sc_hs__clkbuf_1
Xoutput28 net28 VGND VGND VPWR VPWR SWN[4] sky130_fd_sc_hs__clkbuf_1
Xoutput39 net39 VGND VGND VPWR VPWR SWP[7] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_13_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_40_ net4 net5 net14 VGND VGND VPWR VPWR net6 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_23_ net15 _08_ _09_ VGND VGND VPWR VPWR _00_ sky130_fd_sc_hs__o21a_1
XPHY_EDGE_ROW_7_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xoutput18 net18 VGND VGND VPWR VPWR DATA[2] sky130_fd_sc_hs__clkbuf_1
Xoutput29 net29 VGND VGND VPWR VPWR SWN[5] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_22_ _07_ net14 net3 VGND VGND VPWR VPWR _09_ sky130_fd_sc_hs__or3b_1
XFILLER_0_15_116 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_16_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
Xoutput19 net19 VGND VGND VPWR VPWR DATA[3] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_3_44 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_14_94 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_13_64 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_21_ net3 _07_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hs__nand2_1
XFILLER_0_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_3_45 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_13_65 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_20_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[2\] clk_div_0.COUNT\[3\] clk_div_0.COUNT\[0\]
+ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hs__or4bb_1
XFILLER_0_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
Xinput1 CMP_N VGND VGND VPWR VPWR net1 sky130_fd_sc_hs__clkbuf_2
XFILLER_0_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_3_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_56 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
Xinput2 CMP_P VGND VGND VPWR VPWR net2 sky130_fd_sc_hs__buf_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_11_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_14_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_57 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
Xinput3 EN VGND VGND VPWR VPWR net3 sky130_fd_sc_hs__clkbuf_8
XPHY_EDGE_ROW_2_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_0_38 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
Xinput4 RDY VGND VGND VPWR VPWR net4 sky130_fd_sc_hs__buf_2
XTAP_TAPCELL_ROW_10_58 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_0_102 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_0_39 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_10_59 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_59_ net5 net2 net14 VGND VGND VPWR VPWR net32 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_14_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_75_ cyclic_flag_0.FINAL net32 net3 VGND VGND VPWR VPWR net16 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_58_ net6 net2 net14 VGND VGND VPWR VPWR net33 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_6_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_1_40 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_74_ cyclic_flag_0.FINAL net33 net3 VGND VGND VPWR VPWR net17 sky130_fd_sc_hs__dfrtp_1
X_57_ net7 net2 net14 VGND VGND VPWR VPWR net34 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_11_60 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_1_41 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_73_ cyclic_flag_0.FINAL net34 net3 VGND VGND VPWR VPWR net18 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_11_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_56_ net8 net2 net14 VGND VGND VPWR VPWR net35 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_11_61 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_39_ net4 net14 net14 VGND VGND VPWR VPWR net5 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_12_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_72_ cyclic_flag_0.FINAL net35 net3 VGND VGND VPWR VPWR net19 sky130_fd_sc_hs__dfrtp_1
X_55_ net9 net2 net14 VGND VGND VPWR VPWR net36 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_7_52 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_38_ clknet_1_1__leaf_CLK _01_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hs__dfxtp_4
XFILLER_0_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_14_49 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_17_72 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_71_ cyclic_flag_0.FINAL net36 net3 VGND VGND VPWR VPWR net20 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_54_ net10 net2 net14 VGND VGND VPWR VPWR net37 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_7_53 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_37_ clknet_1_1__leaf_CLK _00_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hs__dfxtp_1
XTAP_TAPCELL_ROW_17_73 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_70_ cyclic_flag_0.FINAL net37 net3 VGND VGND VPWR VPWR net21 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hs__clkbuf_16
X_53_ net11 net2 net14 VGND VGND VPWR VPWR net38 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_36_ clk_div_0.COUNT\[3\] _16_ _17_ _10_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hs__o211a_1
X_19_ _06_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_17_74 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_52_ net12 net2 net14 VGND VGND VPWR VPWR net39 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_35_ clk_div_0.COUNT\[3\] _16_ VGND VGND VPWR VPWR _17_ sky130_fd_sc_hs__nand2_1
X_18_ net14 cyclic_flag_0.FINAL VGND VGND VPWR VPWR _06_ sky130_fd_sc_hs__and2_1
XTAP_TAPCELL_ROW_17_75 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_9_102 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_116 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_51_ clknet_1_1__leaf_CLK _05_ VGND VGND VPWR VPWR clk_div_0.COUNT\[3\] sky130_fd_sc_hs__dfxtp_1
X_34_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _16_ sky130_fd_sc_hs__and3_1
XFILLER_0_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_4_46 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_29 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_14_66 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_17_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_50_ clknet_1_0__leaf_CLK _04_ VGND VGND VPWR VPWR clk_div_0.COUNT\[2\] sky130_fd_sc_hs__dfxtp_1
XFILLER_0_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_33_ _15_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hs__clkbuf_1
XFILLER_0_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_5_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_4_47 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_14_67 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_32_ _10_ _14_ VGND VGND VPWR VPWR _15_ sky130_fd_sc_hs__and2_1
XFILLER_0_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_31_ clk_div_0.COUNT\[2\] _12_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hs__xor2_1
XFILLER_0_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_12_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_30_ _08_ _12_ _13_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hs__nor3_1
XFILLER_0_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_9_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_4_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_10 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_12_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_2_42 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_62 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_69_ cyclic_flag_0.FINAL net38 net3 VGND VGND VPWR VPWR net22 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_16_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_2_43 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_12_63 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_68_ cyclic_flag_0.FINAL net39 net3 VGND VGND VPWR VPWR net23 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_4_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput5 net5 VGND VGND VPWR VPWR CF[0] sky130_fd_sc_hs__clkbuf_1
Xclkbuf_1_0__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_0__leaf_CLK sky130_fd_sc_hs__clkbuf_16
XTAP_TAPCELL_ROW_8_54 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_67_ net5 net1 net14 VGND VGND VPWR VPWR net24 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
Xoutput30 net30 VGND VGND VPWR VPWR SWN[6] sky130_fd_sc_hs__clkbuf_1
Xoutput6 net6 VGND VGND VPWR VPWR CF[1] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
.ends

