magic
tech sky130A
magscale 1 2
timestamp 1746016723
<< error_p >>
rect -29 441 29 447
rect -29 407 -17 441
rect -29 401 29 407
rect -29 229 29 235
rect -29 195 -17 229
rect -29 189 29 195
rect -29 17 29 23
rect -29 -17 -17 17
rect -29 -23 29 -17
rect -29 -195 29 -189
rect -29 -229 -17 -195
rect -29 -235 29 -229
rect -29 -407 29 -401
rect -29 -441 -17 -407
rect -29 -447 29 -441
<< nwell >>
rect -109 -460 109 460
<< pmos >>
rect -15 276 15 360
rect -15 64 15 148
rect -15 -148 15 -64
rect -15 -360 15 -276
<< pdiff >>
rect -73 348 -15 360
rect -73 288 -61 348
rect -27 288 -15 348
rect -73 276 -15 288
rect 15 348 73 360
rect 15 288 27 348
rect 61 288 73 348
rect 15 276 73 288
rect -73 136 -15 148
rect -73 76 -61 136
rect -27 76 -15 136
rect -73 64 -15 76
rect 15 136 73 148
rect 15 76 27 136
rect 61 76 73 136
rect 15 64 73 76
rect -73 -76 -15 -64
rect -73 -136 -61 -76
rect -27 -136 -15 -76
rect -73 -148 -15 -136
rect 15 -76 73 -64
rect 15 -136 27 -76
rect 61 -136 73 -76
rect 15 -148 73 -136
rect -73 -288 -15 -276
rect -73 -348 -61 -288
rect -27 -348 -15 -288
rect -73 -360 -15 -348
rect 15 -288 73 -276
rect 15 -348 27 -288
rect 61 -348 73 -288
rect 15 -360 73 -348
<< pdiffc >>
rect -61 288 -27 348
rect 27 288 61 348
rect -61 76 -27 136
rect 27 76 61 136
rect -61 -136 -27 -76
rect 27 -136 61 -76
rect -61 -348 -27 -288
rect 27 -348 61 -288
<< poly >>
rect -33 441 33 457
rect -33 407 -17 441
rect 17 407 33 441
rect -33 391 33 407
rect -15 360 15 391
rect -15 245 15 276
rect -33 229 33 245
rect -33 195 -17 229
rect 17 195 33 229
rect -33 179 33 195
rect -15 148 15 179
rect -15 33 15 64
rect -33 17 33 33
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -33 33 -17
rect -15 -64 15 -33
rect -15 -179 15 -148
rect -33 -195 33 -179
rect -33 -229 -17 -195
rect 17 -229 33 -195
rect -33 -245 33 -229
rect -15 -276 15 -245
rect -15 -391 15 -360
rect -33 -407 33 -391
rect -33 -441 -17 -407
rect 17 -441 33 -407
rect -33 -457 33 -441
<< polycont >>
rect -17 407 17 441
rect -17 195 17 229
rect -17 -17 17 17
rect -17 -229 17 -195
rect -17 -441 17 -407
<< locali >>
rect -33 407 -17 441
rect 17 407 33 441
rect -61 348 -27 364
rect -61 272 -27 288
rect 27 348 61 364
rect 27 272 61 288
rect -33 195 -17 229
rect 17 195 33 229
rect -61 136 -27 152
rect -61 60 -27 76
rect 27 136 61 152
rect 27 60 61 76
rect -33 -17 -17 17
rect 17 -17 33 17
rect -61 -76 -27 -60
rect -61 -152 -27 -136
rect 27 -76 61 -60
rect 27 -152 61 -136
rect -33 -229 -17 -195
rect 17 -229 33 -195
rect -61 -288 -27 -272
rect -61 -364 -27 -348
rect 27 -288 61 -272
rect 27 -364 61 -348
rect -33 -441 -17 -407
rect 17 -441 33 -407
<< viali >>
rect -17 407 17 441
rect -61 288 -27 348
rect 27 288 61 348
rect -17 195 17 229
rect -61 76 -27 136
rect 27 76 61 136
rect -17 -17 17 17
rect -61 -136 -27 -76
rect 27 -136 61 -76
rect -17 -229 17 -195
rect -61 -348 -27 -288
rect 27 -348 61 -288
rect -17 -441 17 -407
<< metal1 >>
rect -29 441 29 447
rect -29 407 -17 441
rect 17 407 29 441
rect -29 401 29 407
rect -67 348 -21 360
rect -67 288 -61 348
rect -27 288 -21 348
rect -67 276 -21 288
rect 21 348 67 360
rect 21 288 27 348
rect 61 288 67 348
rect 21 276 67 288
rect -29 229 29 235
rect -29 195 -17 229
rect 17 195 29 229
rect -29 189 29 195
rect -67 136 -21 148
rect -67 76 -61 136
rect -27 76 -21 136
rect -67 64 -21 76
rect 21 136 67 148
rect 21 76 27 136
rect 61 76 67 136
rect 21 64 67 76
rect -29 17 29 23
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -23 29 -17
rect -67 -76 -21 -64
rect -67 -136 -61 -76
rect -27 -136 -21 -76
rect -67 -148 -21 -136
rect 21 -76 67 -64
rect 21 -136 27 -76
rect 61 -136 67 -76
rect 21 -148 67 -136
rect -29 -195 29 -189
rect -29 -229 -17 -195
rect 17 -229 29 -195
rect -29 -235 29 -229
rect -67 -288 -21 -276
rect -67 -348 -61 -288
rect -27 -348 -21 -288
rect -67 -360 -21 -348
rect 21 -288 67 -276
rect 21 -348 27 -288
rect 61 -348 67 -288
rect 21 -360 67 -348
rect -29 -407 29 -401
rect -29 -441 -17 -407
rect 17 -441 29 -407
rect -29 -447 29 -441
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 4 nf 1 diffcov 100 polycov 20 guard 0 glc 0 grc 1 gtc 0 gbc 0 tbcov 20 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
