magic
tech sky130A
magscale 1 2
timestamp 1746016723
<< error_p >>
rect -29 603 29 609
rect -29 569 -17 603
rect -29 563 29 569
rect -29 391 29 397
rect -29 357 -17 391
rect -29 351 29 357
rect -29 283 29 289
rect -29 249 -17 283
rect -29 243 29 249
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -249 29 -243
rect -29 -283 -17 -249
rect -29 -289 29 -283
rect -29 -357 29 -351
rect -29 -391 -17 -357
rect -29 -397 29 -391
rect -29 -569 29 -563
rect -29 -603 -17 -569
rect -29 -609 29 -603
<< nwell >>
rect -211 -741 211 741
<< pmos >>
rect -15 438 15 522
rect -15 118 15 202
rect -15 -202 15 -118
rect -15 -522 15 -438
<< pdiff >>
rect -73 510 -15 522
rect -73 450 -61 510
rect -27 450 -15 510
rect -73 438 -15 450
rect 15 510 73 522
rect 15 450 27 510
rect 61 450 73 510
rect 15 438 73 450
rect -73 190 -15 202
rect -73 130 -61 190
rect -27 130 -15 190
rect -73 118 -15 130
rect 15 190 73 202
rect 15 130 27 190
rect 61 130 73 190
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -190 -61 -130
rect -27 -190 -15 -130
rect -73 -202 -15 -190
rect 15 -130 73 -118
rect 15 -190 27 -130
rect 61 -190 73 -130
rect 15 -202 73 -190
rect -73 -450 -15 -438
rect -73 -510 -61 -450
rect -27 -510 -15 -450
rect -73 -522 -15 -510
rect 15 -450 73 -438
rect 15 -510 27 -450
rect 61 -510 73 -450
rect 15 -522 73 -510
<< pdiffc >>
rect -61 450 -27 510
rect 27 450 61 510
rect -61 130 -27 190
rect 27 130 61 190
rect -61 -190 -27 -130
rect 27 -190 61 -130
rect -61 -510 -27 -450
rect 27 -510 61 -450
<< nsubdiff >>
rect -175 671 -79 705
rect 79 671 175 705
rect -175 609 -141 671
rect 141 609 175 671
rect -175 -671 -141 -609
rect 141 -671 175 -609
rect -175 -705 -79 -671
rect 79 -705 175 -671
<< nsubdiffcont >>
rect -79 671 79 705
rect -175 -609 -141 609
rect 141 -609 175 609
rect -79 -705 79 -671
<< poly >>
rect -33 603 33 619
rect -33 569 -17 603
rect 17 569 33 603
rect -33 553 33 569
rect -15 522 15 553
rect -15 407 15 438
rect -33 391 33 407
rect -33 357 -17 391
rect 17 357 33 391
rect -33 341 33 357
rect -33 283 33 299
rect -33 249 -17 283
rect 17 249 33 283
rect -33 233 33 249
rect -15 202 15 233
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -233 15 -202
rect -33 -249 33 -233
rect -33 -283 -17 -249
rect 17 -283 33 -249
rect -33 -299 33 -283
rect -33 -357 33 -341
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -33 -407 33 -391
rect -15 -438 15 -407
rect -15 -553 15 -522
rect -33 -569 33 -553
rect -33 -603 -17 -569
rect 17 -603 33 -569
rect -33 -619 33 -603
<< polycont >>
rect -17 569 17 603
rect -17 357 17 391
rect -17 249 17 283
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -283 17 -249
rect -17 -391 17 -357
rect -17 -603 17 -569
<< locali >>
rect -175 671 -79 705
rect 79 671 175 705
rect -175 609 -141 671
rect 141 609 175 671
rect -33 569 -17 603
rect 17 569 33 603
rect -61 510 -27 526
rect -61 434 -27 450
rect 27 510 61 526
rect 27 434 61 450
rect -33 357 -17 391
rect 17 357 33 391
rect -33 249 -17 283
rect 17 249 33 283
rect -61 190 -27 206
rect -61 114 -27 130
rect 27 190 61 206
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -206 -27 -190
rect 27 -130 61 -114
rect 27 -206 61 -190
rect -33 -283 -17 -249
rect 17 -283 33 -249
rect -33 -391 -17 -357
rect 17 -391 33 -357
rect -61 -450 -27 -434
rect -61 -526 -27 -510
rect 27 -450 61 -434
rect 27 -526 61 -510
rect -33 -603 -17 -569
rect 17 -603 33 -569
rect -175 -671 -141 -609
rect 141 -671 175 -609
rect -175 -705 -79 -671
rect 79 -705 175 -671
<< viali >>
rect -17 569 17 603
rect -61 450 -27 510
rect 27 450 61 510
rect -17 357 17 391
rect -17 249 17 283
rect -61 130 -27 190
rect 27 130 61 190
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -190 -27 -130
rect 27 -190 61 -130
rect -17 -283 17 -249
rect -17 -391 17 -357
rect -61 -510 -27 -450
rect 27 -510 61 -450
rect -17 -603 17 -569
<< metal1 >>
rect -29 603 29 609
rect -29 569 -17 603
rect 17 569 29 603
rect -29 563 29 569
rect -67 510 -21 522
rect -67 450 -61 510
rect -27 450 -21 510
rect -67 438 -21 450
rect 21 510 67 522
rect 21 450 27 510
rect 61 450 67 510
rect 21 438 67 450
rect -29 391 29 397
rect -29 357 -17 391
rect 17 357 29 391
rect -29 351 29 357
rect -29 283 29 289
rect -29 249 -17 283
rect 17 249 29 283
rect -29 243 29 249
rect -67 190 -21 202
rect -67 130 -61 190
rect -27 130 -21 190
rect -67 118 -21 130
rect 21 190 67 202
rect 21 130 27 190
rect 61 130 67 190
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -190 -61 -130
rect -27 -190 -21 -130
rect -67 -202 -21 -190
rect 21 -130 67 -118
rect 21 -190 27 -130
rect 61 -190 67 -130
rect 21 -202 67 -190
rect -29 -249 29 -243
rect -29 -283 -17 -249
rect 17 -283 29 -249
rect -29 -289 29 -283
rect -29 -357 29 -351
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -397 29 -391
rect -67 -450 -21 -438
rect -67 -510 -61 -450
rect -27 -510 -21 -450
rect -67 -522 -21 -510
rect 21 -450 67 -438
rect 21 -510 27 -450
rect 61 -510 67 -450
rect 21 -522 67 -510
rect -29 -569 29 -563
rect -29 -603 -17 -569
rect 17 -603 29 -569
rect -29 -609 29 -603
<< properties >>
string FIXED_BBOX -158 -688 158 688
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 4 nf 1 diffcov 100 polycov 20 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
