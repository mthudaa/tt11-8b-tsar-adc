magic
tech sky130A
magscale 1 2
timestamp 1746020920
<< nwell >>
rect -246 -4389 246 4389
<< pmos >>
rect -50 3870 50 4170
rect -50 3334 50 3634
rect -50 2798 50 3098
rect -50 2262 50 2562
rect -50 1726 50 2026
rect -50 1190 50 1490
rect -50 654 50 954
rect -50 118 50 418
rect -50 -418 50 -118
rect -50 -954 50 -654
rect -50 -1490 50 -1190
rect -50 -2026 50 -1726
rect -50 -2562 50 -2262
rect -50 -3098 50 -2798
rect -50 -3634 50 -3334
rect -50 -4170 50 -3870
<< pdiff >>
rect -108 4158 -50 4170
rect -108 3882 -96 4158
rect -62 3882 -50 4158
rect -108 3870 -50 3882
rect 50 4158 108 4170
rect 50 3882 62 4158
rect 96 3882 108 4158
rect 50 3870 108 3882
rect -108 3622 -50 3634
rect -108 3346 -96 3622
rect -62 3346 -50 3622
rect -108 3334 -50 3346
rect 50 3622 108 3634
rect 50 3346 62 3622
rect 96 3346 108 3622
rect 50 3334 108 3346
rect -108 3086 -50 3098
rect -108 2810 -96 3086
rect -62 2810 -50 3086
rect -108 2798 -50 2810
rect 50 3086 108 3098
rect 50 2810 62 3086
rect 96 2810 108 3086
rect 50 2798 108 2810
rect -108 2550 -50 2562
rect -108 2274 -96 2550
rect -62 2274 -50 2550
rect -108 2262 -50 2274
rect 50 2550 108 2562
rect 50 2274 62 2550
rect 96 2274 108 2550
rect 50 2262 108 2274
rect -108 2014 -50 2026
rect -108 1738 -96 2014
rect -62 1738 -50 2014
rect -108 1726 -50 1738
rect 50 2014 108 2026
rect 50 1738 62 2014
rect 96 1738 108 2014
rect 50 1726 108 1738
rect -108 1478 -50 1490
rect -108 1202 -96 1478
rect -62 1202 -50 1478
rect -108 1190 -50 1202
rect 50 1478 108 1490
rect 50 1202 62 1478
rect 96 1202 108 1478
rect 50 1190 108 1202
rect -108 942 -50 954
rect -108 666 -96 942
rect -62 666 -50 942
rect -108 654 -50 666
rect 50 942 108 954
rect 50 666 62 942
rect 96 666 108 942
rect 50 654 108 666
rect -108 406 -50 418
rect -108 130 -96 406
rect -62 130 -50 406
rect -108 118 -50 130
rect 50 406 108 418
rect 50 130 62 406
rect 96 130 108 406
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -406 -96 -130
rect -62 -406 -50 -130
rect -108 -418 -50 -406
rect 50 -130 108 -118
rect 50 -406 62 -130
rect 96 -406 108 -130
rect 50 -418 108 -406
rect -108 -666 -50 -654
rect -108 -942 -96 -666
rect -62 -942 -50 -666
rect -108 -954 -50 -942
rect 50 -666 108 -654
rect 50 -942 62 -666
rect 96 -942 108 -666
rect 50 -954 108 -942
rect -108 -1202 -50 -1190
rect -108 -1478 -96 -1202
rect -62 -1478 -50 -1202
rect -108 -1490 -50 -1478
rect 50 -1202 108 -1190
rect 50 -1478 62 -1202
rect 96 -1478 108 -1202
rect 50 -1490 108 -1478
rect -108 -1738 -50 -1726
rect -108 -2014 -96 -1738
rect -62 -2014 -50 -1738
rect -108 -2026 -50 -2014
rect 50 -1738 108 -1726
rect 50 -2014 62 -1738
rect 96 -2014 108 -1738
rect 50 -2026 108 -2014
rect -108 -2274 -50 -2262
rect -108 -2550 -96 -2274
rect -62 -2550 -50 -2274
rect -108 -2562 -50 -2550
rect 50 -2274 108 -2262
rect 50 -2550 62 -2274
rect 96 -2550 108 -2274
rect 50 -2562 108 -2550
rect -108 -2810 -50 -2798
rect -108 -3086 -96 -2810
rect -62 -3086 -50 -2810
rect -108 -3098 -50 -3086
rect 50 -2810 108 -2798
rect 50 -3086 62 -2810
rect 96 -3086 108 -2810
rect 50 -3098 108 -3086
rect -108 -3346 -50 -3334
rect -108 -3622 -96 -3346
rect -62 -3622 -50 -3346
rect -108 -3634 -50 -3622
rect 50 -3346 108 -3334
rect 50 -3622 62 -3346
rect 96 -3622 108 -3346
rect 50 -3634 108 -3622
rect -108 -3882 -50 -3870
rect -108 -4158 -96 -3882
rect -62 -4158 -50 -3882
rect -108 -4170 -50 -4158
rect 50 -3882 108 -3870
rect 50 -4158 62 -3882
rect 96 -4158 108 -3882
rect 50 -4170 108 -4158
<< pdiffc >>
rect -96 3882 -62 4158
rect 62 3882 96 4158
rect -96 3346 -62 3622
rect 62 3346 96 3622
rect -96 2810 -62 3086
rect 62 2810 96 3086
rect -96 2274 -62 2550
rect 62 2274 96 2550
rect -96 1738 -62 2014
rect 62 1738 96 2014
rect -96 1202 -62 1478
rect 62 1202 96 1478
rect -96 666 -62 942
rect 62 666 96 942
rect -96 130 -62 406
rect 62 130 96 406
rect -96 -406 -62 -130
rect 62 -406 96 -130
rect -96 -942 -62 -666
rect 62 -942 96 -666
rect -96 -1478 -62 -1202
rect 62 -1478 96 -1202
rect -96 -2014 -62 -1738
rect 62 -2014 96 -1738
rect -96 -2550 -62 -2274
rect 62 -2550 96 -2274
rect -96 -3086 -62 -2810
rect 62 -3086 96 -2810
rect -96 -3622 -62 -3346
rect 62 -3622 96 -3346
rect -96 -4158 -62 -3882
rect 62 -4158 96 -3882
<< nsubdiff >>
rect -210 4319 -114 4353
rect 114 4319 210 4353
rect -210 4257 -176 4319
rect 176 4257 210 4319
rect -210 -4319 -176 -4257
rect 176 -4319 210 -4257
rect -210 -4353 -114 -4319
rect 114 -4353 210 -4319
<< nsubdiffcont >>
rect -114 4319 114 4353
rect -210 -4257 -176 4257
rect 176 -4257 210 4257
rect -114 -4353 114 -4319
<< poly >>
rect -50 4251 50 4267
rect -50 4217 -34 4251
rect 34 4217 50 4251
rect -50 4170 50 4217
rect -50 3823 50 3870
rect -50 3789 -34 3823
rect 34 3789 50 3823
rect -50 3773 50 3789
rect -50 3715 50 3731
rect -50 3681 -34 3715
rect 34 3681 50 3715
rect -50 3634 50 3681
rect -50 3287 50 3334
rect -50 3253 -34 3287
rect 34 3253 50 3287
rect -50 3237 50 3253
rect -50 3179 50 3195
rect -50 3145 -34 3179
rect 34 3145 50 3179
rect -50 3098 50 3145
rect -50 2751 50 2798
rect -50 2717 -34 2751
rect 34 2717 50 2751
rect -50 2701 50 2717
rect -50 2643 50 2659
rect -50 2609 -34 2643
rect 34 2609 50 2643
rect -50 2562 50 2609
rect -50 2215 50 2262
rect -50 2181 -34 2215
rect 34 2181 50 2215
rect -50 2165 50 2181
rect -50 2107 50 2123
rect -50 2073 -34 2107
rect 34 2073 50 2107
rect -50 2026 50 2073
rect -50 1679 50 1726
rect -50 1645 -34 1679
rect 34 1645 50 1679
rect -50 1629 50 1645
rect -50 1571 50 1587
rect -50 1537 -34 1571
rect 34 1537 50 1571
rect -50 1490 50 1537
rect -50 1143 50 1190
rect -50 1109 -34 1143
rect 34 1109 50 1143
rect -50 1093 50 1109
rect -50 1035 50 1051
rect -50 1001 -34 1035
rect 34 1001 50 1035
rect -50 954 50 1001
rect -50 607 50 654
rect -50 573 -34 607
rect 34 573 50 607
rect -50 557 50 573
rect -50 499 50 515
rect -50 465 -34 499
rect 34 465 50 499
rect -50 418 50 465
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -465 50 -418
rect -50 -499 -34 -465
rect 34 -499 50 -465
rect -50 -515 50 -499
rect -50 -573 50 -557
rect -50 -607 -34 -573
rect 34 -607 50 -573
rect -50 -654 50 -607
rect -50 -1001 50 -954
rect -50 -1035 -34 -1001
rect 34 -1035 50 -1001
rect -50 -1051 50 -1035
rect -50 -1109 50 -1093
rect -50 -1143 -34 -1109
rect 34 -1143 50 -1109
rect -50 -1190 50 -1143
rect -50 -1537 50 -1490
rect -50 -1571 -34 -1537
rect 34 -1571 50 -1537
rect -50 -1587 50 -1571
rect -50 -1645 50 -1629
rect -50 -1679 -34 -1645
rect 34 -1679 50 -1645
rect -50 -1726 50 -1679
rect -50 -2073 50 -2026
rect -50 -2107 -34 -2073
rect 34 -2107 50 -2073
rect -50 -2123 50 -2107
rect -50 -2181 50 -2165
rect -50 -2215 -34 -2181
rect 34 -2215 50 -2181
rect -50 -2262 50 -2215
rect -50 -2609 50 -2562
rect -50 -2643 -34 -2609
rect 34 -2643 50 -2609
rect -50 -2659 50 -2643
rect -50 -2717 50 -2701
rect -50 -2751 -34 -2717
rect 34 -2751 50 -2717
rect -50 -2798 50 -2751
rect -50 -3145 50 -3098
rect -50 -3179 -34 -3145
rect 34 -3179 50 -3145
rect -50 -3195 50 -3179
rect -50 -3253 50 -3237
rect -50 -3287 -34 -3253
rect 34 -3287 50 -3253
rect -50 -3334 50 -3287
rect -50 -3681 50 -3634
rect -50 -3715 -34 -3681
rect 34 -3715 50 -3681
rect -50 -3731 50 -3715
rect -50 -3789 50 -3773
rect -50 -3823 -34 -3789
rect 34 -3823 50 -3789
rect -50 -3870 50 -3823
rect -50 -4217 50 -4170
rect -50 -4251 -34 -4217
rect 34 -4251 50 -4217
rect -50 -4267 50 -4251
<< polycont >>
rect -34 4217 34 4251
rect -34 3789 34 3823
rect -34 3681 34 3715
rect -34 3253 34 3287
rect -34 3145 34 3179
rect -34 2717 34 2751
rect -34 2609 34 2643
rect -34 2181 34 2215
rect -34 2073 34 2107
rect -34 1645 34 1679
rect -34 1537 34 1571
rect -34 1109 34 1143
rect -34 1001 34 1035
rect -34 573 34 607
rect -34 465 34 499
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -499 34 -465
rect -34 -607 34 -573
rect -34 -1035 34 -1001
rect -34 -1143 34 -1109
rect -34 -1571 34 -1537
rect -34 -1679 34 -1645
rect -34 -2107 34 -2073
rect -34 -2215 34 -2181
rect -34 -2643 34 -2609
rect -34 -2751 34 -2717
rect -34 -3179 34 -3145
rect -34 -3287 34 -3253
rect -34 -3715 34 -3681
rect -34 -3823 34 -3789
rect -34 -4251 34 -4217
<< locali >>
rect -210 4319 -114 4353
rect 114 4319 210 4353
rect -210 4257 -176 4319
rect 176 4257 210 4319
rect -50 4217 -34 4251
rect 34 4217 50 4251
rect -96 4158 -62 4174
rect -96 3866 -62 3882
rect 62 4158 96 4174
rect 62 3866 96 3882
rect -50 3789 -34 3823
rect 34 3789 50 3823
rect -50 3681 -34 3715
rect 34 3681 50 3715
rect -96 3622 -62 3638
rect -96 3330 -62 3346
rect 62 3622 96 3638
rect 62 3330 96 3346
rect -50 3253 -34 3287
rect 34 3253 50 3287
rect -50 3145 -34 3179
rect 34 3145 50 3179
rect -96 3086 -62 3102
rect -96 2794 -62 2810
rect 62 3086 96 3102
rect 62 2794 96 2810
rect -50 2717 -34 2751
rect 34 2717 50 2751
rect -50 2609 -34 2643
rect 34 2609 50 2643
rect -96 2550 -62 2566
rect -96 2258 -62 2274
rect 62 2550 96 2566
rect 62 2258 96 2274
rect -50 2181 -34 2215
rect 34 2181 50 2215
rect -50 2073 -34 2107
rect 34 2073 50 2107
rect -96 2014 -62 2030
rect -96 1722 -62 1738
rect 62 2014 96 2030
rect 62 1722 96 1738
rect -50 1645 -34 1679
rect 34 1645 50 1679
rect -50 1537 -34 1571
rect 34 1537 50 1571
rect -96 1478 -62 1494
rect -96 1186 -62 1202
rect 62 1478 96 1494
rect 62 1186 96 1202
rect -50 1109 -34 1143
rect 34 1109 50 1143
rect -50 1001 -34 1035
rect 34 1001 50 1035
rect -96 942 -62 958
rect -96 650 -62 666
rect 62 942 96 958
rect 62 650 96 666
rect -50 573 -34 607
rect 34 573 50 607
rect -50 465 -34 499
rect 34 465 50 499
rect -96 406 -62 422
rect -96 114 -62 130
rect 62 406 96 422
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -422 -62 -406
rect 62 -130 96 -114
rect 62 -422 96 -406
rect -50 -499 -34 -465
rect 34 -499 50 -465
rect -50 -607 -34 -573
rect 34 -607 50 -573
rect -96 -666 -62 -650
rect -96 -958 -62 -942
rect 62 -666 96 -650
rect 62 -958 96 -942
rect -50 -1035 -34 -1001
rect 34 -1035 50 -1001
rect -50 -1143 -34 -1109
rect 34 -1143 50 -1109
rect -96 -1202 -62 -1186
rect -96 -1494 -62 -1478
rect 62 -1202 96 -1186
rect 62 -1494 96 -1478
rect -50 -1571 -34 -1537
rect 34 -1571 50 -1537
rect -50 -1679 -34 -1645
rect 34 -1679 50 -1645
rect -96 -1738 -62 -1722
rect -96 -2030 -62 -2014
rect 62 -1738 96 -1722
rect 62 -2030 96 -2014
rect -50 -2107 -34 -2073
rect 34 -2107 50 -2073
rect -50 -2215 -34 -2181
rect 34 -2215 50 -2181
rect -96 -2274 -62 -2258
rect -96 -2566 -62 -2550
rect 62 -2274 96 -2258
rect 62 -2566 96 -2550
rect -50 -2643 -34 -2609
rect 34 -2643 50 -2609
rect -50 -2751 -34 -2717
rect 34 -2751 50 -2717
rect -96 -2810 -62 -2794
rect -96 -3102 -62 -3086
rect 62 -2810 96 -2794
rect 62 -3102 96 -3086
rect -50 -3179 -34 -3145
rect 34 -3179 50 -3145
rect -50 -3287 -34 -3253
rect 34 -3287 50 -3253
rect -96 -3346 -62 -3330
rect -96 -3638 -62 -3622
rect 62 -3346 96 -3330
rect 62 -3638 96 -3622
rect -50 -3715 -34 -3681
rect 34 -3715 50 -3681
rect -50 -3823 -34 -3789
rect 34 -3823 50 -3789
rect -96 -3882 -62 -3866
rect -96 -4174 -62 -4158
rect 62 -3882 96 -3866
rect 62 -4174 96 -4158
rect -50 -4251 -34 -4217
rect 34 -4251 50 -4217
rect -210 -4319 -176 -4257
rect 176 -4319 210 -4257
rect -210 -4353 -114 -4319
rect 114 -4353 210 -4319
<< viali >>
rect -34 4217 34 4251
rect -96 3882 -62 4158
rect 62 3882 96 4158
rect -34 3789 34 3823
rect -34 3681 34 3715
rect -96 3346 -62 3622
rect 62 3346 96 3622
rect -34 3253 34 3287
rect -34 3145 34 3179
rect -96 2810 -62 3086
rect 62 2810 96 3086
rect -34 2717 34 2751
rect -34 2609 34 2643
rect -96 2274 -62 2550
rect 62 2274 96 2550
rect -34 2181 34 2215
rect -34 2073 34 2107
rect -96 1738 -62 2014
rect 62 1738 96 2014
rect -34 1645 34 1679
rect -34 1537 34 1571
rect -96 1202 -62 1478
rect 62 1202 96 1478
rect -34 1109 34 1143
rect -34 1001 34 1035
rect -96 666 -62 942
rect 62 666 96 942
rect -34 573 34 607
rect -34 465 34 499
rect -96 130 -62 406
rect 62 130 96 406
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -406 -62 -130
rect 62 -406 96 -130
rect -34 -499 34 -465
rect -34 -607 34 -573
rect -96 -942 -62 -666
rect 62 -942 96 -666
rect -34 -1035 34 -1001
rect -34 -1143 34 -1109
rect -96 -1478 -62 -1202
rect 62 -1478 96 -1202
rect -34 -1571 34 -1537
rect -34 -1679 34 -1645
rect -96 -2014 -62 -1738
rect 62 -2014 96 -1738
rect -34 -2107 34 -2073
rect -34 -2215 34 -2181
rect -96 -2550 -62 -2274
rect 62 -2550 96 -2274
rect -34 -2643 34 -2609
rect -34 -2751 34 -2717
rect -96 -3086 -62 -2810
rect 62 -3086 96 -2810
rect -34 -3179 34 -3145
rect -34 -3287 34 -3253
rect -96 -3622 -62 -3346
rect 62 -3622 96 -3346
rect -34 -3715 34 -3681
rect -34 -3823 34 -3789
rect -96 -4158 -62 -3882
rect 62 -4158 96 -3882
rect -34 -4251 34 -4217
<< metal1 >>
rect -46 4251 46 4257
rect -46 4217 -34 4251
rect 34 4217 46 4251
rect -46 4211 46 4217
rect -102 4158 -56 4170
rect -102 3882 -96 4158
rect -62 3882 -56 4158
rect -102 3870 -56 3882
rect 56 4158 102 4170
rect 56 3882 62 4158
rect 96 3882 102 4158
rect 56 3870 102 3882
rect -46 3823 46 3829
rect -46 3789 -34 3823
rect 34 3789 46 3823
rect -46 3783 46 3789
rect -46 3715 46 3721
rect -46 3681 -34 3715
rect 34 3681 46 3715
rect -46 3675 46 3681
rect -102 3622 -56 3634
rect -102 3346 -96 3622
rect -62 3346 -56 3622
rect -102 3334 -56 3346
rect 56 3622 102 3634
rect 56 3346 62 3622
rect 96 3346 102 3622
rect 56 3334 102 3346
rect -46 3287 46 3293
rect -46 3253 -34 3287
rect 34 3253 46 3287
rect -46 3247 46 3253
rect -46 3179 46 3185
rect -46 3145 -34 3179
rect 34 3145 46 3179
rect -46 3139 46 3145
rect -102 3086 -56 3098
rect -102 2810 -96 3086
rect -62 2810 -56 3086
rect -102 2798 -56 2810
rect 56 3086 102 3098
rect 56 2810 62 3086
rect 96 2810 102 3086
rect 56 2798 102 2810
rect -46 2751 46 2757
rect -46 2717 -34 2751
rect 34 2717 46 2751
rect -46 2711 46 2717
rect -46 2643 46 2649
rect -46 2609 -34 2643
rect 34 2609 46 2643
rect -46 2603 46 2609
rect -102 2550 -56 2562
rect -102 2274 -96 2550
rect -62 2274 -56 2550
rect -102 2262 -56 2274
rect 56 2550 102 2562
rect 56 2274 62 2550
rect 96 2274 102 2550
rect 56 2262 102 2274
rect -46 2215 46 2221
rect -46 2181 -34 2215
rect 34 2181 46 2215
rect -46 2175 46 2181
rect -46 2107 46 2113
rect -46 2073 -34 2107
rect 34 2073 46 2107
rect -46 2067 46 2073
rect -102 2014 -56 2026
rect -102 1738 -96 2014
rect -62 1738 -56 2014
rect -102 1726 -56 1738
rect 56 2014 102 2026
rect 56 1738 62 2014
rect 96 1738 102 2014
rect 56 1726 102 1738
rect -46 1679 46 1685
rect -46 1645 -34 1679
rect 34 1645 46 1679
rect -46 1639 46 1645
rect -46 1571 46 1577
rect -46 1537 -34 1571
rect 34 1537 46 1571
rect -46 1531 46 1537
rect -102 1478 -56 1490
rect -102 1202 -96 1478
rect -62 1202 -56 1478
rect -102 1190 -56 1202
rect 56 1478 102 1490
rect 56 1202 62 1478
rect 96 1202 102 1478
rect 56 1190 102 1202
rect -46 1143 46 1149
rect -46 1109 -34 1143
rect 34 1109 46 1143
rect -46 1103 46 1109
rect -46 1035 46 1041
rect -46 1001 -34 1035
rect 34 1001 46 1035
rect -46 995 46 1001
rect -102 942 -56 954
rect -102 666 -96 942
rect -62 666 -56 942
rect -102 654 -56 666
rect 56 942 102 954
rect 56 666 62 942
rect 96 666 102 942
rect 56 654 102 666
rect -46 607 46 613
rect -46 573 -34 607
rect 34 573 46 607
rect -46 567 46 573
rect -46 499 46 505
rect -46 465 -34 499
rect 34 465 46 499
rect -46 459 46 465
rect -102 406 -56 418
rect -102 130 -96 406
rect -62 130 -56 406
rect -102 118 -56 130
rect 56 406 102 418
rect 56 130 62 406
rect 96 130 102 406
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -406 -96 -130
rect -62 -406 -56 -130
rect -102 -418 -56 -406
rect 56 -130 102 -118
rect 56 -406 62 -130
rect 96 -406 102 -130
rect 56 -418 102 -406
rect -46 -465 46 -459
rect -46 -499 -34 -465
rect 34 -499 46 -465
rect -46 -505 46 -499
rect -46 -573 46 -567
rect -46 -607 -34 -573
rect 34 -607 46 -573
rect -46 -613 46 -607
rect -102 -666 -56 -654
rect -102 -942 -96 -666
rect -62 -942 -56 -666
rect -102 -954 -56 -942
rect 56 -666 102 -654
rect 56 -942 62 -666
rect 96 -942 102 -666
rect 56 -954 102 -942
rect -46 -1001 46 -995
rect -46 -1035 -34 -1001
rect 34 -1035 46 -1001
rect -46 -1041 46 -1035
rect -46 -1109 46 -1103
rect -46 -1143 -34 -1109
rect 34 -1143 46 -1109
rect -46 -1149 46 -1143
rect -102 -1202 -56 -1190
rect -102 -1478 -96 -1202
rect -62 -1478 -56 -1202
rect -102 -1490 -56 -1478
rect 56 -1202 102 -1190
rect 56 -1478 62 -1202
rect 96 -1478 102 -1202
rect 56 -1490 102 -1478
rect -46 -1537 46 -1531
rect -46 -1571 -34 -1537
rect 34 -1571 46 -1537
rect -46 -1577 46 -1571
rect -46 -1645 46 -1639
rect -46 -1679 -34 -1645
rect 34 -1679 46 -1645
rect -46 -1685 46 -1679
rect -102 -1738 -56 -1726
rect -102 -2014 -96 -1738
rect -62 -2014 -56 -1738
rect -102 -2026 -56 -2014
rect 56 -1738 102 -1726
rect 56 -2014 62 -1738
rect 96 -2014 102 -1738
rect 56 -2026 102 -2014
rect -46 -2073 46 -2067
rect -46 -2107 -34 -2073
rect 34 -2107 46 -2073
rect -46 -2113 46 -2107
rect -46 -2181 46 -2175
rect -46 -2215 -34 -2181
rect 34 -2215 46 -2181
rect -46 -2221 46 -2215
rect -102 -2274 -56 -2262
rect -102 -2550 -96 -2274
rect -62 -2550 -56 -2274
rect -102 -2562 -56 -2550
rect 56 -2274 102 -2262
rect 56 -2550 62 -2274
rect 96 -2550 102 -2274
rect 56 -2562 102 -2550
rect -46 -2609 46 -2603
rect -46 -2643 -34 -2609
rect 34 -2643 46 -2609
rect -46 -2649 46 -2643
rect -46 -2717 46 -2711
rect -46 -2751 -34 -2717
rect 34 -2751 46 -2717
rect -46 -2757 46 -2751
rect -102 -2810 -56 -2798
rect -102 -3086 -96 -2810
rect -62 -3086 -56 -2810
rect -102 -3098 -56 -3086
rect 56 -2810 102 -2798
rect 56 -3086 62 -2810
rect 96 -3086 102 -2810
rect 56 -3098 102 -3086
rect -46 -3145 46 -3139
rect -46 -3179 -34 -3145
rect 34 -3179 46 -3145
rect -46 -3185 46 -3179
rect -46 -3253 46 -3247
rect -46 -3287 -34 -3253
rect 34 -3287 46 -3253
rect -46 -3293 46 -3287
rect -102 -3346 -56 -3334
rect -102 -3622 -96 -3346
rect -62 -3622 -56 -3346
rect -102 -3634 -56 -3622
rect 56 -3346 102 -3334
rect 56 -3622 62 -3346
rect 96 -3622 102 -3346
rect 56 -3634 102 -3622
rect -46 -3681 46 -3675
rect -46 -3715 -34 -3681
rect 34 -3715 46 -3681
rect -46 -3721 46 -3715
rect -46 -3789 46 -3783
rect -46 -3823 -34 -3789
rect 34 -3823 46 -3789
rect -46 -3829 46 -3823
rect -102 -3882 -56 -3870
rect -102 -4158 -96 -3882
rect -62 -4158 -56 -3882
rect -102 -4170 -56 -4158
rect 56 -3882 102 -3870
rect 56 -4158 62 -3882
rect 96 -4158 102 -3882
rect 56 -4170 102 -4158
rect -46 -4217 46 -4211
rect -46 -4251 -34 -4217
rect 34 -4251 46 -4217
rect -46 -4257 46 -4251
<< properties >>
string FIXED_BBOX -193 -4336 193 4336
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.5 m 16 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
